magic
tech sky130A
magscale 1 2
timestamp 1624002729
<< nwell >>
rect -66 7703 5538 8577
rect -66 6075 5538 6949
rect -66 4447 5538 5321
rect -66 2819 5538 3693
rect -66 1191 5538 2065
<< locali >>
rect 1759 8585 1892 8719
rect 1037 7636 1081 7713
rect 1325 7636 1369 7713
rect 1613 7636 1657 7713
rect 1901 7636 1945 7713
rect 2189 7636 2233 7713
rect 2477 7636 2521 7713
rect 2765 7636 2809 7713
rect 3053 7636 3097 7713
rect 3341 7636 3385 7713
rect 3629 7636 3673 7713
rect 3871 7642 4001 7676
rect 1037 6939 1081 7016
rect 1325 6939 1369 7016
rect 1613 6939 1657 7016
rect 1901 6939 1945 7016
rect 2189 6939 2233 7016
rect 2477 6939 2521 7016
rect 2765 6939 2809 7016
rect 3053 6939 3097 7016
rect 3341 6939 3385 7016
rect 3629 6939 3673 7016
rect 3871 6976 4001 7010
rect 991 5311 1121 5388
rect 1279 5311 1409 5388
rect 1567 5311 1697 5388
rect 1855 5311 1985 5388
rect 2143 5311 2273 5388
rect 2431 5311 2561 5388
rect 2719 5311 2849 5388
rect 3007 5311 3137 5388
rect 3295 5311 3425 5388
rect 3583 5311 3713 5388
rect 3871 5348 4001 5382
rect 991 4380 1121 4457
rect 1279 4380 1409 4457
rect 1567 4380 1697 4457
rect 1855 4380 1985 4457
rect 2143 4380 2273 4457
rect 2431 4380 2561 4457
rect 2719 4380 2849 4457
rect 3007 4380 3137 4457
rect 3295 4380 3425 4457
rect 3583 4380 3713 4457
rect 3871 4386 4001 4420
rect 1364 2158 1627 2207
rect 2335 2092 2465 2200
rect 3002 2018 3142 2087
rect 1753 1124 1895 1201
rect 2046 1130 2193 1164
<< viali >>
rect 2047 8752 2081 8786
rect 1183 8678 1217 8712
rect 1087 8604 1121 8638
rect 2431 8604 2465 8638
rect 2527 8604 2561 8638
rect 2815 8604 2849 8638
rect 3391 8604 3425 8638
rect 3583 8604 3617 8638
rect 4255 8604 4289 8638
rect 127 8530 161 8564
rect 895 8530 929 8564
rect 2719 8530 2753 8564
rect 893 7641 933 7681
rect 4543 7642 4577 7676
rect 800 6976 834 7010
rect 4543 6976 4577 7010
rect 127 6014 161 6048
rect 895 6014 929 6048
rect 1087 6014 1121 6048
rect 1759 6014 1793 6048
rect 2431 6014 2465 6048
rect 2527 6014 2561 6048
rect 2815 6014 2849 6048
rect 3391 6014 3425 6048
rect 3583 6014 3617 6048
rect 4159 6014 4193 6048
rect 1180 5933 1220 5973
rect 1951 5940 1985 5974
rect 2143 5940 2177 5974
rect 2719 5940 2753 5974
rect 797 5345 837 5385
rect 4543 5348 4577 5382
rect 799 4386 833 4420
rect 4543 4386 4577 4420
rect 2527 3868 2561 3902
rect 2911 3794 2945 3828
rect 3295 3794 3329 3828
rect 3967 3794 4001 3828
rect 2335 3720 2369 3754
rect 3295 3720 3329 3754
rect 3103 3646 3137 3680
rect 127 3424 161 3458
rect 3775 2980 3809 3014
rect 2911 2832 2945 2866
rect 4231 2832 4265 2866
rect 391 2758 425 2792
rect 2431 2758 2465 2792
rect 2719 2758 2753 2792
rect 3103 2758 3137 2792
rect 2623 2684 2657 2718
rect 3103 2684 3137 2718
rect 127 2610 161 2644
rect 127 2240 161 2274
rect 991 2240 1025 2274
rect 2047 2240 2081 2274
rect 2623 2240 2657 2274
rect 487 2166 521 2200
rect 799 2166 833 2200
rect 1759 2166 1793 2200
rect 2143 2092 2177 2126
rect 3487 2092 3521 2126
rect 3967 2092 4001 2126
rect 3391 2018 3425 2052
rect 3775 2018 3809 2052
rect 3871 2018 3905 2052
rect 3487 1870 3521 1904
rect 4231 1796 4265 1830
rect 1759 1352 1793 1386
rect 127 1204 161 1238
rect 895 1204 929 1238
rect 487 1130 521 1164
rect 1087 1130 1121 1164
rect 2815 1130 2849 1164
rect 1087 1056 1121 1090
rect 3007 1056 3041 1090
<< metal1 >>
rect 0 8954 5472 8977
rect 0 8876 149 8954
rect 610 8876 5472 8954
rect 0 8829 5472 8876
rect 785 8744 791 8796
rect 843 8792 849 8796
rect 843 8786 2093 8792
rect 843 8752 2047 8786
rect 2081 8752 2093 8786
rect 843 8746 2093 8752
rect 843 8744 849 8746
rect 1171 8712 1275 8718
rect 1171 8678 1183 8712
rect 1217 8678 1275 8712
rect 1171 8672 1275 8678
rect 1011 8638 1133 8644
rect 1229 8642 1275 8672
rect 3437 8672 5495 8718
rect 3437 8644 3483 8672
rect 1011 8604 1087 8638
rect 1121 8604 1133 8638
rect 1011 8598 1133 8604
rect -23 8564 941 8570
rect -23 8530 127 8564
rect 161 8530 895 8564
rect 929 8530 941 8564
rect -23 8524 941 8530
rect 887 8426 939 8432
rect 1011 8423 1057 8598
rect 1220 8590 1226 8642
rect 1278 8590 1284 8642
rect 2419 8638 2861 8644
rect 2419 8604 2431 8638
rect 2465 8604 2527 8638
rect 2561 8604 2815 8638
rect 2849 8604 2861 8638
rect 2419 8598 2861 8604
rect 3379 8638 3483 8644
rect 3379 8604 3391 8638
rect 3425 8604 3483 8638
rect 3379 8598 3483 8604
rect 3533 8638 3629 8644
rect 3533 8604 3583 8638
rect 3617 8604 3629 8638
rect 3533 8598 3629 8604
rect 4243 8638 5495 8644
rect 4243 8604 4255 8638
rect 4289 8604 5495 8638
rect 4243 8598 5495 8604
rect 1229 8506 1275 8590
rect 3533 8570 3579 8598
rect 2707 8564 3579 8570
rect 2707 8530 2719 8564
rect 2753 8530 3579 8564
rect 2707 8524 3579 8530
rect 939 8377 1057 8423
rect 887 8368 939 8374
rect 0 8209 5472 8265
rect 0 8071 4845 8209
rect 5306 8071 5472 8209
rect 0 8015 5472 8071
rect 1220 7930 1226 7982
rect 1278 7978 1284 7982
rect 1278 7932 4642 7978
rect 1278 7930 1284 7932
rect 881 7635 887 7687
rect 939 7635 945 7687
rect 4596 7682 4642 7932
rect 4531 7676 4644 7682
rect 4531 7642 4543 7676
rect 4577 7642 4644 7676
rect 4531 7636 4644 7642
rect 0 7404 5472 7451
rect 0 7248 149 7404
rect 610 7248 5472 7404
rect 0 7201 5472 7248
rect 881 7115 887 7167
rect 939 7164 945 7167
rect 939 7118 4648 7164
rect 939 7115 945 7118
rect 791 7103 843 7109
rect 791 7045 843 7051
rect 794 7010 840 7045
rect 4602 7016 4648 7118
rect 794 6976 800 7010
rect 834 6976 840 7010
rect 794 6720 840 6976
rect 4531 7010 4648 7016
rect 4531 6976 4543 7010
rect 4577 6976 4648 7010
rect 4531 6970 4648 6976
rect 4059 6720 4065 6723
rect 794 6674 4065 6720
rect 4059 6671 4065 6674
rect 4117 6671 4123 6723
rect 0 6581 5472 6637
rect 0 6443 4845 6581
rect 5306 6443 5472 6581
rect 0 6387 5472 6443
rect 912 6302 918 6354
rect 970 6351 976 6354
rect 970 6305 1692 6351
rect 970 6302 976 6305
rect -23 6048 941 6054
rect -23 6014 127 6048
rect 161 6014 895 6048
rect 929 6014 941 6048
rect -23 6008 941 6014
rect 1010 6048 1133 6054
rect 1010 6014 1087 6048
rect 1121 6014 1133 6048
rect 1010 6008 1133 6014
rect 785 5859 791 5911
rect 843 5908 849 5911
rect 1010 5908 1056 6008
rect 1646 5980 1692 6305
rect 3461 6082 5495 6128
rect 3461 6054 3507 6082
rect 1747 6048 2140 6054
rect 1747 6014 1759 6048
rect 1793 6014 2140 6048
rect 1747 6008 2140 6014
rect 2419 6048 2861 6054
rect 2419 6014 2431 6048
rect 2465 6014 2527 6048
rect 2561 6014 2815 6048
rect 2849 6014 2861 6048
rect 2419 6008 2861 6014
rect 3379 6048 3507 6054
rect 3379 6014 3391 6048
rect 3425 6014 3507 6048
rect 3379 6008 3507 6014
rect 3550 6048 3629 6054
rect 3550 6014 3583 6048
rect 3617 6014 3629 6048
rect 3550 6008 3629 6014
rect 4147 6048 5495 6054
rect 4147 6014 4159 6048
rect 4193 6014 5495 6048
rect 4147 6008 5495 6014
rect 2094 5980 2140 6008
rect 3550 5980 3596 6008
rect 1168 5927 1174 5979
rect 1226 5927 1232 5979
rect 1646 5974 1997 5980
rect 1646 5940 1951 5974
rect 1985 5940 1997 5974
rect 1646 5934 1997 5940
rect 2094 5974 2189 5980
rect 2094 5940 2143 5974
rect 2177 5940 2189 5974
rect 2094 5934 2189 5940
rect 2707 5974 3596 5980
rect 2707 5940 2719 5974
rect 2753 5940 3596 5974
rect 2707 5934 3596 5940
rect 843 5862 1056 5908
rect 843 5859 849 5862
rect 0 5776 5472 5823
rect 0 5620 149 5776
rect 610 5620 5472 5776
rect 0 5573 5472 5620
rect 1174 5539 1226 5545
rect 1226 5490 4635 5536
rect 1174 5481 1226 5487
rect 785 5339 791 5391
rect 843 5339 849 5391
rect 4589 5388 4635 5490
rect 4531 5382 4635 5388
rect 4531 5348 4543 5382
rect 4577 5348 4635 5382
rect 4531 5342 4635 5348
rect 0 4953 5472 5009
rect 0 4815 4845 4953
rect 5306 4815 5472 4953
rect 0 4759 5472 4815
rect 785 4673 791 4725
rect 843 4722 849 4725
rect 843 4676 4620 4722
rect 843 4673 849 4676
rect 794 4426 840 4428
rect 4574 4426 4620 4676
rect 787 4420 845 4426
rect 787 4386 799 4420
rect 833 4386 845 4420
rect 787 4380 845 4386
rect 4531 4420 4620 4426
rect 4531 4386 4543 4420
rect 4577 4386 4620 4420
rect 4531 4380 4620 4386
rect 794 4278 840 4380
rect 918 4311 970 4317
rect 794 4259 918 4278
rect 3828 4278 3834 4281
rect 970 4259 3834 4278
rect 794 4232 3834 4259
rect 3828 4229 3834 4232
rect 3886 4229 3892 4281
rect 0 4148 5472 4195
rect 0 3992 149 4148
rect 610 3992 5472 4148
rect 0 3945 5472 3992
rect 2515 3902 3684 3908
rect 2515 3868 2527 3902
rect 2561 3895 3684 3902
rect 2561 3868 3626 3895
rect 2515 3862 3626 3868
rect 3620 3843 3626 3862
rect 3678 3843 3684 3895
rect 4059 3834 4065 3837
rect 2899 3828 3341 3834
rect 2899 3794 2911 3828
rect 2945 3794 3295 3828
rect 3329 3794 3341 3828
rect 2899 3788 3341 3794
rect 3955 3828 4065 3834
rect 3955 3794 3967 3828
rect 4001 3794 4065 3828
rect 3955 3788 4065 3794
rect 4059 3785 4065 3788
rect 4117 3785 4123 3837
rect 2304 3711 2310 3763
rect 2362 3760 2368 3763
rect 2362 3754 2381 3760
rect 2369 3720 2381 3754
rect 2362 3714 2381 3720
rect 3234 3754 3341 3760
rect 3234 3720 3295 3754
rect 3329 3720 3341 3754
rect 3234 3714 3341 3720
rect 2362 3711 2368 3714
rect 3039 3680 3149 3686
rect 3039 3646 3103 3680
rect 3137 3646 3149 3680
rect 3039 3640 3149 3646
rect 2872 3616 2924 3622
rect 3039 3613 3085 3640
rect 2924 3567 3085 3613
rect 3039 3566 3085 3567
rect 2872 3558 2924 3564
rect 3234 3464 3280 3714
rect -23 3458 3280 3464
rect -23 3424 127 3458
rect 161 3424 3280 3458
rect -23 3418 3280 3424
rect 0 3325 5472 3381
rect 0 3187 4845 3325
rect 5306 3187 5472 3325
rect 0 3131 5472 3187
rect 2872 3041 2924 3047
rect -23 2989 2872 3020
rect 3828 3020 3834 3023
rect -23 2983 2924 2989
rect 3763 3014 3834 3020
rect -23 2974 2921 2983
rect 3763 2980 3775 3014
rect 3809 2980 3834 3014
rect 3763 2974 3834 2980
rect 2195 2900 2846 2946
rect 2195 2798 2241 2900
rect 0 2792 2241 2798
rect 0 2758 391 2792
rect 425 2758 2241 2792
rect 2313 2826 2706 2872
rect 2313 2777 2359 2826
rect 2660 2798 2706 2826
rect 2800 2798 2846 2900
rect 2875 2872 2921 2974
rect 3828 2971 3834 2974
rect 3886 2971 3892 3023
rect 2875 2866 4277 2872
rect 2875 2832 2911 2866
rect 2945 2832 4231 2866
rect 4265 2832 4277 2866
rect 2875 2826 4277 2832
rect 2419 2792 2527 2798
rect 0 2752 2241 2758
rect 2310 2771 2362 2777
rect 2419 2758 2431 2792
rect 2465 2758 2527 2792
rect 2419 2752 2527 2758
rect 2660 2792 2765 2798
rect 2660 2758 2719 2792
rect 2753 2758 2765 2792
rect 2660 2752 2765 2758
rect 2800 2792 3149 2798
rect 2800 2758 3103 2792
rect 3137 2758 3149 2792
rect 2800 2752 3149 2758
rect 2310 2713 2362 2719
rect 2313 2650 2359 2713
rect 0 2644 2359 2650
rect 0 2610 127 2644
rect 161 2610 2359 2644
rect 0 2604 2359 2610
rect 2481 2650 2527 2752
rect 2611 2718 3149 2724
rect 2611 2684 2623 2718
rect 2657 2684 3103 2718
rect 3137 2684 3149 2718
rect 2611 2678 3149 2684
rect 3282 2650 3288 2653
rect 2481 2604 3288 2650
rect 3282 2601 3288 2604
rect 3340 2601 3346 2653
rect 0 2520 5472 2567
rect 0 2364 149 2520
rect 610 2364 5472 2520
rect 0 2317 5472 2364
rect -23 2274 1037 2280
rect -23 2240 127 2274
rect 161 2240 991 2274
rect 1025 2240 1037 2274
rect -23 2234 1037 2240
rect 2035 2274 2669 2280
rect 2035 2240 2047 2274
rect 2081 2240 2623 2274
rect 2657 2240 2669 2274
rect 2035 2234 2669 2240
rect -23 2200 845 2206
rect -23 2166 487 2200
rect 521 2166 799 2200
rect 833 2166 845 2200
rect -23 2160 845 2166
rect 1670 2200 1805 2206
rect 1670 2166 1759 2200
rect 1793 2166 1805 2200
rect 1670 2160 1805 2166
rect 3626 2165 3678 2171
rect 1670 2132 1716 2160
rect -23 2086 1716 2132
rect 1670 1836 1716 2086
rect 2058 2083 2064 2135
rect 2116 2132 2122 2135
rect 2116 2126 2975 2132
rect 2116 2092 2143 2126
rect 2177 2092 2975 2126
rect 2116 2086 2975 2092
rect 2116 2083 2122 2086
rect 2929 1984 2975 2086
rect 3282 2083 3288 2135
rect 3340 2132 3346 2135
rect 3340 2126 3567 2132
rect 3340 2092 3487 2126
rect 3521 2092 3567 2126
rect 3678 2126 4050 2132
rect 3678 2113 3967 2126
rect 3626 2107 3967 2113
rect 3340 2086 3567 2092
rect 3629 2092 3967 2107
rect 4001 2092 4050 2126
rect 3629 2086 4050 2092
rect 3340 2083 3346 2086
rect 3629 2058 3675 2086
rect 3379 2052 3675 2058
rect 3379 2018 3391 2052
rect 3425 2018 3675 2052
rect 3379 2012 3675 2018
rect 3719 2052 3821 2058
rect 3719 2018 3775 2052
rect 3809 2018 3821 2052
rect 3719 2012 3821 2018
rect 3859 2052 3917 2058
rect 3859 2018 3871 2052
rect 3905 2018 3917 2052
rect 3955 2037 4001 2086
rect 3859 2012 3917 2018
rect 3719 1984 3765 2012
rect 2929 1945 3765 1984
rect 2930 1938 3765 1945
rect 3859 1910 3905 2012
rect 3475 1904 3905 1910
rect 3475 1870 3487 1904
rect 3521 1878 3905 1904
rect 3521 1870 3904 1878
rect 3475 1864 3904 1870
rect 1670 1830 4277 1836
rect 1670 1796 4231 1830
rect 4265 1796 4277 1830
rect 1670 1790 4277 1796
rect 0 1697 5472 1753
rect 0 1559 4845 1697
rect 5306 1559 5472 1697
rect 0 1503 5472 1559
rect 2058 1392 2064 1395
rect 1747 1386 2064 1392
rect 1747 1352 1759 1386
rect 1793 1352 2064 1386
rect 1747 1346 2064 1352
rect 2058 1343 2064 1346
rect 2116 1343 2122 1395
rect -23 1238 941 1244
rect -23 1204 127 1238
rect 161 1204 895 1238
rect 929 1204 941 1238
rect -23 1198 941 1204
rect -23 1164 1133 1170
rect -23 1130 487 1164
rect 521 1130 1087 1164
rect 1121 1130 1133 1164
rect -23 1124 1133 1130
rect 2803 1164 5495 1170
rect 2803 1130 2815 1164
rect 2849 1130 5495 1164
rect 2803 1124 5495 1130
rect -23 1090 3058 1096
rect -23 1056 1087 1090
rect 1121 1056 3007 1090
rect 3041 1056 3058 1090
rect -23 1050 3058 1056
rect 0 892 5472 939
rect 0 831 127 892
rect 641 831 5472 892
rect 0 791 5472 831
<< via1 >>
rect 149 8876 610 8954
rect 791 8744 843 8796
rect 887 8374 939 8426
rect 1226 8590 1278 8642
rect 4845 8071 5306 8209
rect 1226 7930 1278 7982
rect 887 7681 939 7687
rect 887 7641 893 7681
rect 893 7641 933 7681
rect 933 7641 939 7681
rect 887 7635 939 7641
rect 149 7248 610 7404
rect 887 7115 939 7167
rect 791 7051 843 7103
rect 4065 6671 4117 6723
rect 4845 6443 5306 6581
rect 918 6302 970 6354
rect 791 5859 843 5911
rect 1174 5973 1226 5979
rect 1174 5933 1180 5973
rect 1180 5933 1220 5973
rect 1220 5933 1226 5973
rect 1174 5927 1226 5933
rect 149 5620 610 5776
rect 1174 5487 1226 5539
rect 791 5385 843 5391
rect 791 5345 797 5385
rect 797 5345 837 5385
rect 837 5345 843 5385
rect 791 5339 843 5345
rect 4845 4815 5306 4953
rect 791 4673 843 4725
rect 918 4259 970 4311
rect 3834 4229 3886 4281
rect 149 3992 610 4148
rect 3626 3843 3678 3895
rect 4065 3785 4117 3837
rect 2310 3754 2362 3763
rect 2310 3720 2335 3754
rect 2335 3720 2362 3754
rect 2310 3711 2362 3720
rect 2872 3564 2924 3616
rect 4845 3187 5306 3325
rect 2872 2989 2924 3041
rect 3834 2971 3886 3023
rect 2310 2719 2362 2771
rect 3288 2601 3340 2653
rect 149 2364 610 2520
rect 2064 2083 2116 2135
rect 3288 2083 3340 2135
rect 3626 2113 3678 2165
rect 4845 1559 5306 1697
rect 2064 1343 2116 1395
rect 127 831 641 892
<< metal2 >>
rect 0 8954 699 8997
rect 0 8876 149 8954
rect 610 8876 699 8954
rect 0 7404 699 8876
rect 791 8796 843 8802
rect 791 8738 843 8744
rect 0 7248 149 7404
rect 610 7248 699 7404
rect 0 5776 699 7248
rect 794 7103 840 8738
rect 1226 8642 1278 8648
rect 1226 8584 1278 8590
rect 881 8374 887 8426
rect 939 8374 945 8426
rect 890 7693 936 8374
rect 1229 7988 1275 8584
rect 4773 8209 5472 8997
rect 4773 8071 4845 8209
rect 5306 8071 5472 8209
rect 1226 7982 1278 7988
rect 1226 7924 1278 7930
rect 887 7687 939 7693
rect 887 7629 939 7635
rect 890 7173 936 7629
rect 887 7167 939 7173
rect 887 7109 939 7115
rect 785 7051 791 7103
rect 843 7051 849 7103
rect 4065 6723 4117 6729
rect 4065 6665 4117 6671
rect 918 6354 970 6360
rect 918 6296 970 6302
rect 791 5911 843 5917
rect 791 5853 843 5859
rect 0 5620 149 5776
rect 610 5620 699 5776
rect 0 4148 699 5620
rect 794 5397 840 5853
rect 791 5391 843 5397
rect 791 5333 843 5339
rect 794 4731 840 5333
rect 791 4725 843 4731
rect 791 4667 843 4673
rect 921 4311 967 6296
rect 1174 5979 1226 5985
rect 1174 5921 1226 5927
rect 1177 5539 1223 5921
rect 1168 5487 1174 5539
rect 1226 5487 1232 5539
rect 912 4259 918 4311
rect 970 4259 976 4311
rect 3834 4281 3886 4287
rect 3834 4223 3886 4229
rect 0 3992 149 4148
rect 610 3992 699 4148
rect 0 2520 699 3992
rect 3626 3895 3678 3901
rect 3626 3837 3678 3843
rect 2310 3763 2362 3769
rect 2310 3705 2362 3711
rect 2313 2771 2359 3705
rect 2866 3564 2872 3616
rect 2924 3564 2930 3616
rect 2875 3041 2921 3564
rect 2866 2989 2872 3041
rect 2924 2989 2930 3041
rect 2304 2719 2310 2771
rect 2362 2719 2368 2771
rect 3288 2653 3340 2659
rect 3288 2595 3340 2601
rect 0 2364 149 2520
rect 610 2364 699 2520
rect 0 892 699 2364
rect 3291 2141 3337 2595
rect 3629 2165 3675 3837
rect 3837 3029 3883 4223
rect 4068 3843 4114 6665
rect 4773 6581 5472 8071
rect 4773 6443 4845 6581
rect 5306 6443 5472 6581
rect 4773 4953 5472 6443
rect 4773 4815 4845 4953
rect 5306 4815 5472 4953
rect 4065 3837 4117 3843
rect 4065 3779 4117 3785
rect 4773 3325 5472 4815
rect 4773 3187 4845 3325
rect 5306 3187 5472 3325
rect 3834 3023 3886 3029
rect 3834 2965 3886 2971
rect 2064 2135 2116 2141
rect 2064 2077 2116 2083
rect 3288 2135 3340 2141
rect 3620 2113 3626 2165
rect 3678 2113 3684 2165
rect 3288 2077 3340 2083
rect 2067 1401 2113 2077
rect 4773 1697 5472 3187
rect 4773 1559 4845 1697
rect 5306 1559 5472 1697
rect 2064 1395 2116 1401
rect 2064 1337 2116 1343
rect 0 831 127 892
rect 641 831 699 892
rect 0 791 699 831
rect 4773 791 5472 1559
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_4 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624002729
transform 1 0 360 0 -1 2442
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_3
timestamp 1624002729
transform 1 0 0 0 -1 2442
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_1
timestamp 1624002729
transform 1 0 360 0 1 814
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0
timestamp 1624002729
transform 1 0 0 0 1 814
box -66 -43 258 897
use sky130_fd_sc_hvl__mux2_1  sky130_fd_sc_hvl__mux2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624002729
transform -1 0 1824 0 1 814
box -66 -43 1122 897
use sky130_fd_sc_hvl__and2_1  sky130_fd_sc_hvl__and2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624002729
transform 1 0 768 0 -1 2442
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  sky130_fd_sc_hvl__or2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624002729
transform 1 0 1440 0 -1 2442
box -66 -43 738 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624002729
transform 1 0 1824 0 1 814
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_1
timestamp 1624002729
transform 1 0 2112 0 -1 2442
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624002729
transform 1 0 2112 0 1 814
box -66 -43 834 897
use sky130_fd_sc_hvl__nor2_1  sky130_fd_sc_hvl__nor2_1_1 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624002729
transform 1 0 3552 0 -1 2442
box -66 -43 546 897
use sky130_fd_sc_hvl__nor2_1  sky130_fd_sc_hvl__nor2_1_0
timestamp 1624002729
transform 1 0 3072 0 -1 2442
box -66 -43 546 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_2
timestamp 1624002729
transform 1 0 2976 0 1 814
box -66 -43 258 897
use sky130_fd_sc_hvl__and2_1  sky130_fd_sc_hvl__and2_1_1
timestamp 1624002729
transform 1 0 2400 0 -1 2442
box -66 -43 738 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_7
timestamp 1624002729
transform 1 0 4200 0 -1 2442
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_3 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624002729
transform 1 0 4704 0 -1 2442
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_1
timestamp 1624002729
transform 1 0 4704 0 1 814
box -66 -43 834 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_6
timestamp 1624002729
transform 1 0 360 0 1 2442
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_5
timestamp 1624002729
transform 1 0 0 0 1 2442
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_5
timestamp 1624002729
transform 1 0 768 0 1 2442
box -66 -43 834 897
use sky130_fd_sc_hvl__nand2_1  sky130_fd_sc_hvl__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1624002729
transform 1 0 2304 0 1 2442
box -66 -43 546 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_6
timestamp 1624002729
transform 1 0 1536 0 1 2442
box -66 -43 834 897
use sky130_fd_sc_hvl__mux2_1  sky130_fd_sc_hvl__mux2_1_1
timestamp 1624002729
transform -1 0 3840 0 1 2442
box -66 -43 1122 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_8
timestamp 1624002729
transform 1 0 4200 0 1 2442
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_7
timestamp 1624002729
transform 1 0 4704 0 1 2442
box -66 -43 834 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_9
timestamp 1624002729
transform 1 0 0 0 -1 4070
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_9
timestamp 1624002729
transform 1 0 768 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  sky130_fd_sc_hvl__and2_1_2
timestamp 1624002729
transform 1 0 2304 0 -1 4070
box -66 -43 738 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_10
timestamp 1624002729
transform 1 0 1536 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__mux2_1  sky130_fd_sc_hvl__mux2_1_2
timestamp 1624002729
transform -1 0 4032 0 -1 4070
box -66 -43 1122 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_11
timestamp 1624002729
transform 1 0 4704 0 -1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_12
timestamp 1624002729
transform 1 0 0 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_2
timestamp 1624002729
transform 1 0 768 0 1 4070
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_3
timestamp 1624002729
transform 1 0 1056 0 1 4070
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_4
timestamp 1624002729
transform 1 0 1344 0 1 4070
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_5
timestamp 1624002729
transform 1 0 1632 0 1 4070
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_6
timestamp 1624002729
transform 1 0 1920 0 1 4070
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_7
timestamp 1624002729
transform 1 0 2208 0 1 4070
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_8
timestamp 1624002729
transform 1 0 2496 0 1 4070
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_9
timestamp 1624002729
transform 1 0 2784 0 1 4070
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_10
timestamp 1624002729
transform 1 0 3072 0 1 4070
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_11
timestamp 1624002729
transform 1 0 3360 0 1 4070
box -66 -43 354 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_13
timestamp 1624002729
transform 1 0 4704 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_12
timestamp 1624002729
transform 1 0 3648 0 1 4070
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_1
timestamp 1624002729
transform 1 0 3936 0 1 4070
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_14
timestamp 1624002729
transform 1 0 0 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_13
timestamp 1624002729
transform 1 0 768 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_14
timestamp 1624002729
transform 1 0 1056 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_15
timestamp 1624002729
transform 1 0 1344 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_16
timestamp 1624002729
transform 1 0 1632 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_17
timestamp 1624002729
transform 1 0 1920 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_18
timestamp 1624002729
transform 1 0 2208 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_19
timestamp 1624002729
transform 1 0 2496 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_20
timestamp 1624002729
transform 1 0 2784 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_21
timestamp 1624002729
transform 1 0 3072 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_22
timestamp 1624002729
transform 1 0 3360 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_15
timestamp 1624002729
transform 1 0 4704 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_23
timestamp 1624002729
transform 1 0 3648 0 -1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_2
timestamp 1624002729
transform 1 0 3936 0 -1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_10
timestamp 1624002729
transform 1 0 0 0 1 5698
box -66 -43 258 897
use sky130_fd_sc_hvl__mux2_1  sky130_fd_sc_hvl__mux2_1_3
timestamp 1624002729
transform -1 0 1824 0 1 5698
box -66 -43 1122 897
use sky130_fd_sc_hvl__or2_1  sky130_fd_sc_hvl__or2_1_1
timestamp 1624002729
transform 1 0 1824 0 1 5698
box -66 -43 738 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_24
timestamp 1624002729
transform 1 0 2496 0 1 5698
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_3
timestamp 1624002729
transform 1 0 2784 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_4
timestamp 1624002729
transform 1 0 3552 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_17
timestamp 1624002729
transform 1 0 4704 0 1 5698
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_20
timestamp 1624002729
transform 1 0 0 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_18
timestamp 1624002729
transform 1 0 0 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_25
timestamp 1624002729
transform 1 0 768 0 -1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_26
timestamp 1624002729
transform 1 0 1056 0 -1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_36
timestamp 1624002729
transform 1 0 768 0 1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_37
timestamp 1624002729
transform 1 0 1056 0 1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_27
timestamp 1624002729
transform 1 0 1344 0 -1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_28
timestamp 1624002729
transform 1 0 1632 0 -1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_29
timestamp 1624002729
transform 1 0 1920 0 -1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_30
timestamp 1624002729
transform 1 0 2208 0 -1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_38
timestamp 1624002729
transform 1 0 1344 0 1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_39
timestamp 1624002729
transform 1 0 1632 0 1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_40
timestamp 1624002729
transform 1 0 1920 0 1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_41
timestamp 1624002729
transform 1 0 2208 0 1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_31
timestamp 1624002729
transform 1 0 2496 0 -1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_32
timestamp 1624002729
transform 1 0 2784 0 -1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_33
timestamp 1624002729
transform 1 0 3072 0 -1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_34
timestamp 1624002729
transform 1 0 3360 0 -1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_42
timestamp 1624002729
transform 1 0 2496 0 1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_43
timestamp 1624002729
transform 1 0 2784 0 1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_44
timestamp 1624002729
transform 1 0 3072 0 1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_45
timestamp 1624002729
transform 1 0 3360 0 1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_21
timestamp 1624002729
transform 1 0 4704 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_19
timestamp 1624002729
transform 1 0 4704 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_35
timestamp 1624002729
transform 1 0 3648 0 -1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_46
timestamp 1624002729
transform 1 0 3648 0 1 7326
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_5
timestamp 1624002729
transform 1 0 3936 0 -1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_6
timestamp 1624002729
transform 1 0 3936 0 1 7326
box -66 -43 834 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_11
timestamp 1624002729
transform 1 0 0 0 -1 8954
box -66 -43 258 897
use sky130_fd_sc_hvl__mux2_1  sky130_fd_sc_hvl__mux2_1_4
timestamp 1624002729
transform -1 0 1824 0 -1 8954
box -66 -43 1122 897
use sky130_fd_sc_hvl__and2_1  sky130_fd_sc_hvl__and2_1_3
timestamp 1624002729
transform 1 0 1824 0 -1 8954
box -66 -43 738 897
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_47
timestamp 1624002729
transform 1 0 2496 0 -1 8954
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_7
timestamp 1624002729
transform 1 0 2784 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_8
timestamp 1624002729
transform 1 0 3552 0 -1 8954
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_23
timestamp 1624002729
transform 1 0 4704 0 -1 8954
box -66 -43 834 897
<< labels >>
flabel metal1 3545 2086 3547 2132 1 FreeSans 400 0 0 0 hs_control
flabel metal1 4041 2086 4043 2132 1 FreeSans 400 0 0 0 ls_control
flabel via1 2098 2086 2100 2132 1 FreeSans 400 0 0 0 timeout
flabel metal1 -23 2160 -21 2206 1 FreeSans 400 0 0 0 overcurrent
port 7 n
flabel metal1 -23 2234 -21 2280 1 FreeSans 400 0 0 0 oc_en
port 6 n
flabel metal1 -23 2086 -21 2132 1 FreeSans 400 0 0 0 cycle_end
port 1 n
flabel metal1 -23 1198 -21 1244 1 FreeSans 400 0 0 0 timeout_sel
port 17 n
flabel metal1 -23 1124 -21 1170 1 FreeSans 400 0 0 0 timeout_int
port 15 n
flabel metal1 -23 1050 -21 1096 1 FreeSans 400 0 0 0 timeout_ext
port 14 n
flabel metal1 5493 1124 5495 1170 1 FreeSans 400 0 0 0 timeout_out
port 16 n
flabel metal1 0 2604 2 2650 1 FreeSans 400 0 0 0 sw_en
port 12 n
flabel metal1 0 2752 2 2798 1 FreeSans 400 0 0 0 pmos_val
port 11 n
flabel metal1 -23 2974 -21 3020 1 FreeSans 400 0 0 0 sw_override
port 13 n
flabel via1 3856 2974 3858 3020 1 FreeSans 400 0 0 0 pmos_dly_in
flabel metal1 -23 3418 -21 3464 1 FreeSans 400 0 0 0 nmos_val
port 5 n
flabel metal1 4023 3788 4024 3834 1 FreeSans 400 0 0 0 nmos_dly_in
flabel metal1 4531 4380 4533 4426 1 FreeSans 400 0 0 0 pmos_dly_m
flabel metal1 -23 6008 -21 6054 1 FreeSans 400 0 0 0 pmos_dt
port 10 n
flabel metal1 5493 6008 5495 6054 1 FreeSans 400 0 0 0 pmos_drv
port 8 n
flabel metal1 5493 6082 5495 6128 1 FreeSans 400 0 0 0 pmos_drv_n
port 9 n
flabel metal1 5493 8598 5495 8644 1 FreeSans 400 0 0 0 nmos_drv
port 2 n
flabel metal1 5493 8672 5495 8718 1 FreeSans 400 0 0 0 nmos_drv_n
port 3 n
flabel metal1 s 0 791 4 939 0 FreeSans 400 0 0 0 vss
port 19 nsew
flabel metal1 s 0 1503 4 1753 0 FreeSans 400 0 0 0 vdd
port 18 nsew
flabel metal1 -23 8524 -21 8570 1 FreeSans 400 0 0 0 nmos_dt
port 4 n
<< end >>
