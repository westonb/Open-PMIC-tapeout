magic
tech sky130A
magscale 1 2
timestamp 1624002729
<< error_p >>
rect -7031 566 7031 600
rect -7061 -566 7061 566
rect -7031 -600 7031 -566
<< nwell >>
rect -7031 -600 7031 600
<< mvpmos >>
rect -6937 -500 -6737 500
rect -6679 -500 -6479 500
rect -6421 -500 -6221 500
rect -6163 -500 -5963 500
rect -5905 -500 -5705 500
rect -5647 -500 -5447 500
rect -5389 -500 -5189 500
rect -5131 -500 -4931 500
rect -4873 -500 -4673 500
rect -4615 -500 -4415 500
rect -4357 -500 -4157 500
rect -4099 -500 -3899 500
rect -3841 -500 -3641 500
rect -3583 -500 -3383 500
rect -3325 -500 -3125 500
rect -3067 -500 -2867 500
rect -2809 -500 -2609 500
rect -2551 -500 -2351 500
rect -2293 -500 -2093 500
rect -2035 -500 -1835 500
rect -1777 -500 -1577 500
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
rect 1577 -500 1777 500
rect 1835 -500 2035 500
rect 2093 -500 2293 500
rect 2351 -500 2551 500
rect 2609 -500 2809 500
rect 2867 -500 3067 500
rect 3125 -500 3325 500
rect 3383 -500 3583 500
rect 3641 -500 3841 500
rect 3899 -500 4099 500
rect 4157 -500 4357 500
rect 4415 -500 4615 500
rect 4673 -500 4873 500
rect 4931 -500 5131 500
rect 5189 -500 5389 500
rect 5447 -500 5647 500
rect 5705 -500 5905 500
rect 5963 -500 6163 500
rect 6221 -500 6421 500
rect 6479 -500 6679 500
rect 6737 -500 6937 500
<< mvpdiff >>
rect -6995 488 -6937 500
rect -6995 -488 -6983 488
rect -6949 -488 -6937 488
rect -6995 -500 -6937 -488
rect -6737 488 -6679 500
rect -6737 -488 -6725 488
rect -6691 -488 -6679 488
rect -6737 -500 -6679 -488
rect -6479 488 -6421 500
rect -6479 -488 -6467 488
rect -6433 -488 -6421 488
rect -6479 -500 -6421 -488
rect -6221 488 -6163 500
rect -6221 -488 -6209 488
rect -6175 -488 -6163 488
rect -6221 -500 -6163 -488
rect -5963 488 -5905 500
rect -5963 -488 -5951 488
rect -5917 -488 -5905 488
rect -5963 -500 -5905 -488
rect -5705 488 -5647 500
rect -5705 -488 -5693 488
rect -5659 -488 -5647 488
rect -5705 -500 -5647 -488
rect -5447 488 -5389 500
rect -5447 -488 -5435 488
rect -5401 -488 -5389 488
rect -5447 -500 -5389 -488
rect -5189 488 -5131 500
rect -5189 -488 -5177 488
rect -5143 -488 -5131 488
rect -5189 -500 -5131 -488
rect -4931 488 -4873 500
rect -4931 -488 -4919 488
rect -4885 -488 -4873 488
rect -4931 -500 -4873 -488
rect -4673 488 -4615 500
rect -4673 -488 -4661 488
rect -4627 -488 -4615 488
rect -4673 -500 -4615 -488
rect -4415 488 -4357 500
rect -4415 -488 -4403 488
rect -4369 -488 -4357 488
rect -4415 -500 -4357 -488
rect -4157 488 -4099 500
rect -4157 -488 -4145 488
rect -4111 -488 -4099 488
rect -4157 -500 -4099 -488
rect -3899 488 -3841 500
rect -3899 -488 -3887 488
rect -3853 -488 -3841 488
rect -3899 -500 -3841 -488
rect -3641 488 -3583 500
rect -3641 -488 -3629 488
rect -3595 -488 -3583 488
rect -3641 -500 -3583 -488
rect -3383 488 -3325 500
rect -3383 -488 -3371 488
rect -3337 -488 -3325 488
rect -3383 -500 -3325 -488
rect -3125 488 -3067 500
rect -3125 -488 -3113 488
rect -3079 -488 -3067 488
rect -3125 -500 -3067 -488
rect -2867 488 -2809 500
rect -2867 -488 -2855 488
rect -2821 -488 -2809 488
rect -2867 -500 -2809 -488
rect -2609 488 -2551 500
rect -2609 -488 -2597 488
rect -2563 -488 -2551 488
rect -2609 -500 -2551 -488
rect -2351 488 -2293 500
rect -2351 -488 -2339 488
rect -2305 -488 -2293 488
rect -2351 -500 -2293 -488
rect -2093 488 -2035 500
rect -2093 -488 -2081 488
rect -2047 -488 -2035 488
rect -2093 -500 -2035 -488
rect -1835 488 -1777 500
rect -1835 -488 -1823 488
rect -1789 -488 -1777 488
rect -1835 -500 -1777 -488
rect -1577 488 -1519 500
rect -1577 -488 -1565 488
rect -1531 -488 -1519 488
rect -1577 -500 -1519 -488
rect -1319 488 -1261 500
rect -1319 -488 -1307 488
rect -1273 -488 -1261 488
rect -1319 -500 -1261 -488
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
rect 1261 488 1319 500
rect 1261 -488 1273 488
rect 1307 -488 1319 488
rect 1261 -500 1319 -488
rect 1519 488 1577 500
rect 1519 -488 1531 488
rect 1565 -488 1577 488
rect 1519 -500 1577 -488
rect 1777 488 1835 500
rect 1777 -488 1789 488
rect 1823 -488 1835 488
rect 1777 -500 1835 -488
rect 2035 488 2093 500
rect 2035 -488 2047 488
rect 2081 -488 2093 488
rect 2035 -500 2093 -488
rect 2293 488 2351 500
rect 2293 -488 2305 488
rect 2339 -488 2351 488
rect 2293 -500 2351 -488
rect 2551 488 2609 500
rect 2551 -488 2563 488
rect 2597 -488 2609 488
rect 2551 -500 2609 -488
rect 2809 488 2867 500
rect 2809 -488 2821 488
rect 2855 -488 2867 488
rect 2809 -500 2867 -488
rect 3067 488 3125 500
rect 3067 -488 3079 488
rect 3113 -488 3125 488
rect 3067 -500 3125 -488
rect 3325 488 3383 500
rect 3325 -488 3337 488
rect 3371 -488 3383 488
rect 3325 -500 3383 -488
rect 3583 488 3641 500
rect 3583 -488 3595 488
rect 3629 -488 3641 488
rect 3583 -500 3641 -488
rect 3841 488 3899 500
rect 3841 -488 3853 488
rect 3887 -488 3899 488
rect 3841 -500 3899 -488
rect 4099 488 4157 500
rect 4099 -488 4111 488
rect 4145 -488 4157 488
rect 4099 -500 4157 -488
rect 4357 488 4415 500
rect 4357 -488 4369 488
rect 4403 -488 4415 488
rect 4357 -500 4415 -488
rect 4615 488 4673 500
rect 4615 -488 4627 488
rect 4661 -488 4673 488
rect 4615 -500 4673 -488
rect 4873 488 4931 500
rect 4873 -488 4885 488
rect 4919 -488 4931 488
rect 4873 -500 4931 -488
rect 5131 488 5189 500
rect 5131 -488 5143 488
rect 5177 -488 5189 488
rect 5131 -500 5189 -488
rect 5389 488 5447 500
rect 5389 -488 5401 488
rect 5435 -488 5447 488
rect 5389 -500 5447 -488
rect 5647 488 5705 500
rect 5647 -488 5659 488
rect 5693 -488 5705 488
rect 5647 -500 5705 -488
rect 5905 488 5963 500
rect 5905 -488 5917 488
rect 5951 -488 5963 488
rect 5905 -500 5963 -488
rect 6163 488 6221 500
rect 6163 -488 6175 488
rect 6209 -488 6221 488
rect 6163 -500 6221 -488
rect 6421 488 6479 500
rect 6421 -488 6433 488
rect 6467 -488 6479 488
rect 6421 -500 6479 -488
rect 6679 488 6737 500
rect 6679 -488 6691 488
rect 6725 -488 6737 488
rect 6679 -500 6737 -488
rect 6937 488 6995 500
rect 6937 -488 6949 488
rect 6983 -488 6995 488
rect 6937 -500 6995 -488
<< mvpdiffc >>
rect -6983 -488 -6949 488
rect -6725 -488 -6691 488
rect -6467 -488 -6433 488
rect -6209 -488 -6175 488
rect -5951 -488 -5917 488
rect -5693 -488 -5659 488
rect -5435 -488 -5401 488
rect -5177 -488 -5143 488
rect -4919 -488 -4885 488
rect -4661 -488 -4627 488
rect -4403 -488 -4369 488
rect -4145 -488 -4111 488
rect -3887 -488 -3853 488
rect -3629 -488 -3595 488
rect -3371 -488 -3337 488
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect 3337 -488 3371 488
rect 3595 -488 3629 488
rect 3853 -488 3887 488
rect 4111 -488 4145 488
rect 4369 -488 4403 488
rect 4627 -488 4661 488
rect 4885 -488 4919 488
rect 5143 -488 5177 488
rect 5401 -488 5435 488
rect 5659 -488 5693 488
rect 5917 -488 5951 488
rect 6175 -488 6209 488
rect 6433 -488 6467 488
rect 6691 -488 6725 488
rect 6949 -488 6983 488
<< poly >>
rect -6903 581 -6771 597
rect -6903 564 -6887 581
rect -6937 547 -6887 564
rect -6787 564 -6771 581
rect -6645 581 -6513 597
rect -6645 564 -6629 581
rect -6787 547 -6737 564
rect -6937 500 -6737 547
rect -6679 547 -6629 564
rect -6529 564 -6513 581
rect -6387 581 -6255 597
rect -6387 564 -6371 581
rect -6529 547 -6479 564
rect -6679 500 -6479 547
rect -6421 547 -6371 564
rect -6271 564 -6255 581
rect -6129 581 -5997 597
rect -6129 564 -6113 581
rect -6271 547 -6221 564
rect -6421 500 -6221 547
rect -6163 547 -6113 564
rect -6013 564 -5997 581
rect -5871 581 -5739 597
rect -5871 564 -5855 581
rect -6013 547 -5963 564
rect -6163 500 -5963 547
rect -5905 547 -5855 564
rect -5755 564 -5739 581
rect -5613 581 -5481 597
rect -5613 564 -5597 581
rect -5755 547 -5705 564
rect -5905 500 -5705 547
rect -5647 547 -5597 564
rect -5497 564 -5481 581
rect -5355 581 -5223 597
rect -5355 564 -5339 581
rect -5497 547 -5447 564
rect -5647 500 -5447 547
rect -5389 547 -5339 564
rect -5239 564 -5223 581
rect -5097 581 -4965 597
rect -5097 564 -5081 581
rect -5239 547 -5189 564
rect -5389 500 -5189 547
rect -5131 547 -5081 564
rect -4981 564 -4965 581
rect -4839 581 -4707 597
rect -4839 564 -4823 581
rect -4981 547 -4931 564
rect -5131 500 -4931 547
rect -4873 547 -4823 564
rect -4723 564 -4707 581
rect -4581 581 -4449 597
rect -4581 564 -4565 581
rect -4723 547 -4673 564
rect -4873 500 -4673 547
rect -4615 547 -4565 564
rect -4465 564 -4449 581
rect -4323 581 -4191 597
rect -4323 564 -4307 581
rect -4465 547 -4415 564
rect -4615 500 -4415 547
rect -4357 547 -4307 564
rect -4207 564 -4191 581
rect -4065 581 -3933 597
rect -4065 564 -4049 581
rect -4207 547 -4157 564
rect -4357 500 -4157 547
rect -4099 547 -4049 564
rect -3949 564 -3933 581
rect -3807 581 -3675 597
rect -3807 564 -3791 581
rect -3949 547 -3899 564
rect -4099 500 -3899 547
rect -3841 547 -3791 564
rect -3691 564 -3675 581
rect -3549 581 -3417 597
rect -3549 564 -3533 581
rect -3691 547 -3641 564
rect -3841 500 -3641 547
rect -3583 547 -3533 564
rect -3433 564 -3417 581
rect -3291 581 -3159 597
rect -3291 564 -3275 581
rect -3433 547 -3383 564
rect -3583 500 -3383 547
rect -3325 547 -3275 564
rect -3175 564 -3159 581
rect -3033 581 -2901 597
rect -3033 564 -3017 581
rect -3175 547 -3125 564
rect -3325 500 -3125 547
rect -3067 547 -3017 564
rect -2917 564 -2901 581
rect -2775 581 -2643 597
rect -2775 564 -2759 581
rect -2917 547 -2867 564
rect -3067 500 -2867 547
rect -2809 547 -2759 564
rect -2659 564 -2643 581
rect -2517 581 -2385 597
rect -2517 564 -2501 581
rect -2659 547 -2609 564
rect -2809 500 -2609 547
rect -2551 547 -2501 564
rect -2401 564 -2385 581
rect -2259 581 -2127 597
rect -2259 564 -2243 581
rect -2401 547 -2351 564
rect -2551 500 -2351 547
rect -2293 547 -2243 564
rect -2143 564 -2127 581
rect -2001 581 -1869 597
rect -2001 564 -1985 581
rect -2143 547 -2093 564
rect -2293 500 -2093 547
rect -2035 547 -1985 564
rect -1885 564 -1869 581
rect -1743 581 -1611 597
rect -1743 564 -1727 581
rect -1885 547 -1835 564
rect -2035 500 -1835 547
rect -1777 547 -1727 564
rect -1627 564 -1611 581
rect -1485 581 -1353 597
rect -1485 564 -1469 581
rect -1627 547 -1577 564
rect -1777 500 -1577 547
rect -1519 547 -1469 564
rect -1369 564 -1353 581
rect -1227 581 -1095 597
rect -1227 564 -1211 581
rect -1369 547 -1319 564
rect -1519 500 -1319 547
rect -1261 547 -1211 564
rect -1111 564 -1095 581
rect -969 581 -837 597
rect -969 564 -953 581
rect -1111 547 -1061 564
rect -1261 500 -1061 547
rect -1003 547 -953 564
rect -853 564 -837 581
rect -711 581 -579 597
rect -711 564 -695 581
rect -853 547 -803 564
rect -1003 500 -803 547
rect -745 547 -695 564
rect -595 564 -579 581
rect -453 581 -321 597
rect -453 564 -437 581
rect -595 547 -545 564
rect -745 500 -545 547
rect -487 547 -437 564
rect -337 564 -321 581
rect -195 581 -63 597
rect -195 564 -179 581
rect -337 547 -287 564
rect -487 500 -287 547
rect -229 547 -179 564
rect -79 564 -63 581
rect 63 581 195 597
rect 63 564 79 581
rect -79 547 -29 564
rect -229 500 -29 547
rect 29 547 79 564
rect 179 564 195 581
rect 321 581 453 597
rect 321 564 337 581
rect 179 547 229 564
rect 29 500 229 547
rect 287 547 337 564
rect 437 564 453 581
rect 579 581 711 597
rect 579 564 595 581
rect 437 547 487 564
rect 287 500 487 547
rect 545 547 595 564
rect 695 564 711 581
rect 837 581 969 597
rect 837 564 853 581
rect 695 547 745 564
rect 545 500 745 547
rect 803 547 853 564
rect 953 564 969 581
rect 1095 581 1227 597
rect 1095 564 1111 581
rect 953 547 1003 564
rect 803 500 1003 547
rect 1061 547 1111 564
rect 1211 564 1227 581
rect 1353 581 1485 597
rect 1353 564 1369 581
rect 1211 547 1261 564
rect 1061 500 1261 547
rect 1319 547 1369 564
rect 1469 564 1485 581
rect 1611 581 1743 597
rect 1611 564 1627 581
rect 1469 547 1519 564
rect 1319 500 1519 547
rect 1577 547 1627 564
rect 1727 564 1743 581
rect 1869 581 2001 597
rect 1869 564 1885 581
rect 1727 547 1777 564
rect 1577 500 1777 547
rect 1835 547 1885 564
rect 1985 564 2001 581
rect 2127 581 2259 597
rect 2127 564 2143 581
rect 1985 547 2035 564
rect 1835 500 2035 547
rect 2093 547 2143 564
rect 2243 564 2259 581
rect 2385 581 2517 597
rect 2385 564 2401 581
rect 2243 547 2293 564
rect 2093 500 2293 547
rect 2351 547 2401 564
rect 2501 564 2517 581
rect 2643 581 2775 597
rect 2643 564 2659 581
rect 2501 547 2551 564
rect 2351 500 2551 547
rect 2609 547 2659 564
rect 2759 564 2775 581
rect 2901 581 3033 597
rect 2901 564 2917 581
rect 2759 547 2809 564
rect 2609 500 2809 547
rect 2867 547 2917 564
rect 3017 564 3033 581
rect 3159 581 3291 597
rect 3159 564 3175 581
rect 3017 547 3067 564
rect 2867 500 3067 547
rect 3125 547 3175 564
rect 3275 564 3291 581
rect 3417 581 3549 597
rect 3417 564 3433 581
rect 3275 547 3325 564
rect 3125 500 3325 547
rect 3383 547 3433 564
rect 3533 564 3549 581
rect 3675 581 3807 597
rect 3675 564 3691 581
rect 3533 547 3583 564
rect 3383 500 3583 547
rect 3641 547 3691 564
rect 3791 564 3807 581
rect 3933 581 4065 597
rect 3933 564 3949 581
rect 3791 547 3841 564
rect 3641 500 3841 547
rect 3899 547 3949 564
rect 4049 564 4065 581
rect 4191 581 4323 597
rect 4191 564 4207 581
rect 4049 547 4099 564
rect 3899 500 4099 547
rect 4157 547 4207 564
rect 4307 564 4323 581
rect 4449 581 4581 597
rect 4449 564 4465 581
rect 4307 547 4357 564
rect 4157 500 4357 547
rect 4415 547 4465 564
rect 4565 564 4581 581
rect 4707 581 4839 597
rect 4707 564 4723 581
rect 4565 547 4615 564
rect 4415 500 4615 547
rect 4673 547 4723 564
rect 4823 564 4839 581
rect 4965 581 5097 597
rect 4965 564 4981 581
rect 4823 547 4873 564
rect 4673 500 4873 547
rect 4931 547 4981 564
rect 5081 564 5097 581
rect 5223 581 5355 597
rect 5223 564 5239 581
rect 5081 547 5131 564
rect 4931 500 5131 547
rect 5189 547 5239 564
rect 5339 564 5355 581
rect 5481 581 5613 597
rect 5481 564 5497 581
rect 5339 547 5389 564
rect 5189 500 5389 547
rect 5447 547 5497 564
rect 5597 564 5613 581
rect 5739 581 5871 597
rect 5739 564 5755 581
rect 5597 547 5647 564
rect 5447 500 5647 547
rect 5705 547 5755 564
rect 5855 564 5871 581
rect 5997 581 6129 597
rect 5997 564 6013 581
rect 5855 547 5905 564
rect 5705 500 5905 547
rect 5963 547 6013 564
rect 6113 564 6129 581
rect 6255 581 6387 597
rect 6255 564 6271 581
rect 6113 547 6163 564
rect 5963 500 6163 547
rect 6221 547 6271 564
rect 6371 564 6387 581
rect 6513 581 6645 597
rect 6513 564 6529 581
rect 6371 547 6421 564
rect 6221 500 6421 547
rect 6479 547 6529 564
rect 6629 564 6645 581
rect 6771 581 6903 597
rect 6771 564 6787 581
rect 6629 547 6679 564
rect 6479 500 6679 547
rect 6737 547 6787 564
rect 6887 564 6903 581
rect 6887 547 6937 564
rect 6737 500 6937 547
rect -6937 -547 -6737 -500
rect -6937 -564 -6887 -547
rect -6903 -581 -6887 -564
rect -6787 -564 -6737 -547
rect -6679 -547 -6479 -500
rect -6679 -564 -6629 -547
rect -6787 -581 -6771 -564
rect -6903 -597 -6771 -581
rect -6645 -581 -6629 -564
rect -6529 -564 -6479 -547
rect -6421 -547 -6221 -500
rect -6421 -564 -6371 -547
rect -6529 -581 -6513 -564
rect -6645 -597 -6513 -581
rect -6387 -581 -6371 -564
rect -6271 -564 -6221 -547
rect -6163 -547 -5963 -500
rect -6163 -564 -6113 -547
rect -6271 -581 -6255 -564
rect -6387 -597 -6255 -581
rect -6129 -581 -6113 -564
rect -6013 -564 -5963 -547
rect -5905 -547 -5705 -500
rect -5905 -564 -5855 -547
rect -6013 -581 -5997 -564
rect -6129 -597 -5997 -581
rect -5871 -581 -5855 -564
rect -5755 -564 -5705 -547
rect -5647 -547 -5447 -500
rect -5647 -564 -5597 -547
rect -5755 -581 -5739 -564
rect -5871 -597 -5739 -581
rect -5613 -581 -5597 -564
rect -5497 -564 -5447 -547
rect -5389 -547 -5189 -500
rect -5389 -564 -5339 -547
rect -5497 -581 -5481 -564
rect -5613 -597 -5481 -581
rect -5355 -581 -5339 -564
rect -5239 -564 -5189 -547
rect -5131 -547 -4931 -500
rect -5131 -564 -5081 -547
rect -5239 -581 -5223 -564
rect -5355 -597 -5223 -581
rect -5097 -581 -5081 -564
rect -4981 -564 -4931 -547
rect -4873 -547 -4673 -500
rect -4873 -564 -4823 -547
rect -4981 -581 -4965 -564
rect -5097 -597 -4965 -581
rect -4839 -581 -4823 -564
rect -4723 -564 -4673 -547
rect -4615 -547 -4415 -500
rect -4615 -564 -4565 -547
rect -4723 -581 -4707 -564
rect -4839 -597 -4707 -581
rect -4581 -581 -4565 -564
rect -4465 -564 -4415 -547
rect -4357 -547 -4157 -500
rect -4357 -564 -4307 -547
rect -4465 -581 -4449 -564
rect -4581 -597 -4449 -581
rect -4323 -581 -4307 -564
rect -4207 -564 -4157 -547
rect -4099 -547 -3899 -500
rect -4099 -564 -4049 -547
rect -4207 -581 -4191 -564
rect -4323 -597 -4191 -581
rect -4065 -581 -4049 -564
rect -3949 -564 -3899 -547
rect -3841 -547 -3641 -500
rect -3841 -564 -3791 -547
rect -3949 -581 -3933 -564
rect -4065 -597 -3933 -581
rect -3807 -581 -3791 -564
rect -3691 -564 -3641 -547
rect -3583 -547 -3383 -500
rect -3583 -564 -3533 -547
rect -3691 -581 -3675 -564
rect -3807 -597 -3675 -581
rect -3549 -581 -3533 -564
rect -3433 -564 -3383 -547
rect -3325 -547 -3125 -500
rect -3325 -564 -3275 -547
rect -3433 -581 -3417 -564
rect -3549 -597 -3417 -581
rect -3291 -581 -3275 -564
rect -3175 -564 -3125 -547
rect -3067 -547 -2867 -500
rect -3067 -564 -3017 -547
rect -3175 -581 -3159 -564
rect -3291 -597 -3159 -581
rect -3033 -581 -3017 -564
rect -2917 -564 -2867 -547
rect -2809 -547 -2609 -500
rect -2809 -564 -2759 -547
rect -2917 -581 -2901 -564
rect -3033 -597 -2901 -581
rect -2775 -581 -2759 -564
rect -2659 -564 -2609 -547
rect -2551 -547 -2351 -500
rect -2551 -564 -2501 -547
rect -2659 -581 -2643 -564
rect -2775 -597 -2643 -581
rect -2517 -581 -2501 -564
rect -2401 -564 -2351 -547
rect -2293 -547 -2093 -500
rect -2293 -564 -2243 -547
rect -2401 -581 -2385 -564
rect -2517 -597 -2385 -581
rect -2259 -581 -2243 -564
rect -2143 -564 -2093 -547
rect -2035 -547 -1835 -500
rect -2035 -564 -1985 -547
rect -2143 -581 -2127 -564
rect -2259 -597 -2127 -581
rect -2001 -581 -1985 -564
rect -1885 -564 -1835 -547
rect -1777 -547 -1577 -500
rect -1777 -564 -1727 -547
rect -1885 -581 -1869 -564
rect -2001 -597 -1869 -581
rect -1743 -581 -1727 -564
rect -1627 -564 -1577 -547
rect -1519 -547 -1319 -500
rect -1519 -564 -1469 -547
rect -1627 -581 -1611 -564
rect -1743 -597 -1611 -581
rect -1485 -581 -1469 -564
rect -1369 -564 -1319 -547
rect -1261 -547 -1061 -500
rect -1261 -564 -1211 -547
rect -1369 -581 -1353 -564
rect -1485 -597 -1353 -581
rect -1227 -581 -1211 -564
rect -1111 -564 -1061 -547
rect -1003 -547 -803 -500
rect -1003 -564 -953 -547
rect -1111 -581 -1095 -564
rect -1227 -597 -1095 -581
rect -969 -581 -953 -564
rect -853 -564 -803 -547
rect -745 -547 -545 -500
rect -745 -564 -695 -547
rect -853 -581 -837 -564
rect -969 -597 -837 -581
rect -711 -581 -695 -564
rect -595 -564 -545 -547
rect -487 -547 -287 -500
rect -487 -564 -437 -547
rect -595 -581 -579 -564
rect -711 -597 -579 -581
rect -453 -581 -437 -564
rect -337 -564 -287 -547
rect -229 -547 -29 -500
rect -229 -564 -179 -547
rect -337 -581 -321 -564
rect -453 -597 -321 -581
rect -195 -581 -179 -564
rect -79 -564 -29 -547
rect 29 -547 229 -500
rect 29 -564 79 -547
rect -79 -581 -63 -564
rect -195 -597 -63 -581
rect 63 -581 79 -564
rect 179 -564 229 -547
rect 287 -547 487 -500
rect 287 -564 337 -547
rect 179 -581 195 -564
rect 63 -597 195 -581
rect 321 -581 337 -564
rect 437 -564 487 -547
rect 545 -547 745 -500
rect 545 -564 595 -547
rect 437 -581 453 -564
rect 321 -597 453 -581
rect 579 -581 595 -564
rect 695 -564 745 -547
rect 803 -547 1003 -500
rect 803 -564 853 -547
rect 695 -581 711 -564
rect 579 -597 711 -581
rect 837 -581 853 -564
rect 953 -564 1003 -547
rect 1061 -547 1261 -500
rect 1061 -564 1111 -547
rect 953 -581 969 -564
rect 837 -597 969 -581
rect 1095 -581 1111 -564
rect 1211 -564 1261 -547
rect 1319 -547 1519 -500
rect 1319 -564 1369 -547
rect 1211 -581 1227 -564
rect 1095 -597 1227 -581
rect 1353 -581 1369 -564
rect 1469 -564 1519 -547
rect 1577 -547 1777 -500
rect 1577 -564 1627 -547
rect 1469 -581 1485 -564
rect 1353 -597 1485 -581
rect 1611 -581 1627 -564
rect 1727 -564 1777 -547
rect 1835 -547 2035 -500
rect 1835 -564 1885 -547
rect 1727 -581 1743 -564
rect 1611 -597 1743 -581
rect 1869 -581 1885 -564
rect 1985 -564 2035 -547
rect 2093 -547 2293 -500
rect 2093 -564 2143 -547
rect 1985 -581 2001 -564
rect 1869 -597 2001 -581
rect 2127 -581 2143 -564
rect 2243 -564 2293 -547
rect 2351 -547 2551 -500
rect 2351 -564 2401 -547
rect 2243 -581 2259 -564
rect 2127 -597 2259 -581
rect 2385 -581 2401 -564
rect 2501 -564 2551 -547
rect 2609 -547 2809 -500
rect 2609 -564 2659 -547
rect 2501 -581 2517 -564
rect 2385 -597 2517 -581
rect 2643 -581 2659 -564
rect 2759 -564 2809 -547
rect 2867 -547 3067 -500
rect 2867 -564 2917 -547
rect 2759 -581 2775 -564
rect 2643 -597 2775 -581
rect 2901 -581 2917 -564
rect 3017 -564 3067 -547
rect 3125 -547 3325 -500
rect 3125 -564 3175 -547
rect 3017 -581 3033 -564
rect 2901 -597 3033 -581
rect 3159 -581 3175 -564
rect 3275 -564 3325 -547
rect 3383 -547 3583 -500
rect 3383 -564 3433 -547
rect 3275 -581 3291 -564
rect 3159 -597 3291 -581
rect 3417 -581 3433 -564
rect 3533 -564 3583 -547
rect 3641 -547 3841 -500
rect 3641 -564 3691 -547
rect 3533 -581 3549 -564
rect 3417 -597 3549 -581
rect 3675 -581 3691 -564
rect 3791 -564 3841 -547
rect 3899 -547 4099 -500
rect 3899 -564 3949 -547
rect 3791 -581 3807 -564
rect 3675 -597 3807 -581
rect 3933 -581 3949 -564
rect 4049 -564 4099 -547
rect 4157 -547 4357 -500
rect 4157 -564 4207 -547
rect 4049 -581 4065 -564
rect 3933 -597 4065 -581
rect 4191 -581 4207 -564
rect 4307 -564 4357 -547
rect 4415 -547 4615 -500
rect 4415 -564 4465 -547
rect 4307 -581 4323 -564
rect 4191 -597 4323 -581
rect 4449 -581 4465 -564
rect 4565 -564 4615 -547
rect 4673 -547 4873 -500
rect 4673 -564 4723 -547
rect 4565 -581 4581 -564
rect 4449 -597 4581 -581
rect 4707 -581 4723 -564
rect 4823 -564 4873 -547
rect 4931 -547 5131 -500
rect 4931 -564 4981 -547
rect 4823 -581 4839 -564
rect 4707 -597 4839 -581
rect 4965 -581 4981 -564
rect 5081 -564 5131 -547
rect 5189 -547 5389 -500
rect 5189 -564 5239 -547
rect 5081 -581 5097 -564
rect 4965 -597 5097 -581
rect 5223 -581 5239 -564
rect 5339 -564 5389 -547
rect 5447 -547 5647 -500
rect 5447 -564 5497 -547
rect 5339 -581 5355 -564
rect 5223 -597 5355 -581
rect 5481 -581 5497 -564
rect 5597 -564 5647 -547
rect 5705 -547 5905 -500
rect 5705 -564 5755 -547
rect 5597 -581 5613 -564
rect 5481 -597 5613 -581
rect 5739 -581 5755 -564
rect 5855 -564 5905 -547
rect 5963 -547 6163 -500
rect 5963 -564 6013 -547
rect 5855 -581 5871 -564
rect 5739 -597 5871 -581
rect 5997 -581 6013 -564
rect 6113 -564 6163 -547
rect 6221 -547 6421 -500
rect 6221 -564 6271 -547
rect 6113 -581 6129 -564
rect 5997 -597 6129 -581
rect 6255 -581 6271 -564
rect 6371 -564 6421 -547
rect 6479 -547 6679 -500
rect 6479 -564 6529 -547
rect 6371 -581 6387 -564
rect 6255 -597 6387 -581
rect 6513 -581 6529 -564
rect 6629 -564 6679 -547
rect 6737 -547 6937 -500
rect 6737 -564 6787 -547
rect 6629 -581 6645 -564
rect 6513 -597 6645 -581
rect 6771 -581 6787 -564
rect 6887 -564 6937 -547
rect 6887 -581 6903 -564
rect 6771 -597 6903 -581
<< polycont >>
rect -6887 547 -6787 581
rect -6629 547 -6529 581
rect -6371 547 -6271 581
rect -6113 547 -6013 581
rect -5855 547 -5755 581
rect -5597 547 -5497 581
rect -5339 547 -5239 581
rect -5081 547 -4981 581
rect -4823 547 -4723 581
rect -4565 547 -4465 581
rect -4307 547 -4207 581
rect -4049 547 -3949 581
rect -3791 547 -3691 581
rect -3533 547 -3433 581
rect -3275 547 -3175 581
rect -3017 547 -2917 581
rect -2759 547 -2659 581
rect -2501 547 -2401 581
rect -2243 547 -2143 581
rect -1985 547 -1885 581
rect -1727 547 -1627 581
rect -1469 547 -1369 581
rect -1211 547 -1111 581
rect -953 547 -853 581
rect -695 547 -595 581
rect -437 547 -337 581
rect -179 547 -79 581
rect 79 547 179 581
rect 337 547 437 581
rect 595 547 695 581
rect 853 547 953 581
rect 1111 547 1211 581
rect 1369 547 1469 581
rect 1627 547 1727 581
rect 1885 547 1985 581
rect 2143 547 2243 581
rect 2401 547 2501 581
rect 2659 547 2759 581
rect 2917 547 3017 581
rect 3175 547 3275 581
rect 3433 547 3533 581
rect 3691 547 3791 581
rect 3949 547 4049 581
rect 4207 547 4307 581
rect 4465 547 4565 581
rect 4723 547 4823 581
rect 4981 547 5081 581
rect 5239 547 5339 581
rect 5497 547 5597 581
rect 5755 547 5855 581
rect 6013 547 6113 581
rect 6271 547 6371 581
rect 6529 547 6629 581
rect 6787 547 6887 581
rect -6887 -581 -6787 -547
rect -6629 -581 -6529 -547
rect -6371 -581 -6271 -547
rect -6113 -581 -6013 -547
rect -5855 -581 -5755 -547
rect -5597 -581 -5497 -547
rect -5339 -581 -5239 -547
rect -5081 -581 -4981 -547
rect -4823 -581 -4723 -547
rect -4565 -581 -4465 -547
rect -4307 -581 -4207 -547
rect -4049 -581 -3949 -547
rect -3791 -581 -3691 -547
rect -3533 -581 -3433 -547
rect -3275 -581 -3175 -547
rect -3017 -581 -2917 -547
rect -2759 -581 -2659 -547
rect -2501 -581 -2401 -547
rect -2243 -581 -2143 -547
rect -1985 -581 -1885 -547
rect -1727 -581 -1627 -547
rect -1469 -581 -1369 -547
rect -1211 -581 -1111 -547
rect -953 -581 -853 -547
rect -695 -581 -595 -547
rect -437 -581 -337 -547
rect -179 -581 -79 -547
rect 79 -581 179 -547
rect 337 -581 437 -547
rect 595 -581 695 -547
rect 853 -581 953 -547
rect 1111 -581 1211 -547
rect 1369 -581 1469 -547
rect 1627 -581 1727 -547
rect 1885 -581 1985 -547
rect 2143 -581 2243 -547
rect 2401 -581 2501 -547
rect 2659 -581 2759 -547
rect 2917 -581 3017 -547
rect 3175 -581 3275 -547
rect 3433 -581 3533 -547
rect 3691 -581 3791 -547
rect 3949 -581 4049 -547
rect 4207 -581 4307 -547
rect 4465 -581 4565 -547
rect 4723 -581 4823 -547
rect 4981 -581 5081 -547
rect 5239 -581 5339 -547
rect 5497 -581 5597 -547
rect 5755 -581 5855 -547
rect 6013 -581 6113 -547
rect 6271 -581 6371 -547
rect 6529 -581 6629 -547
rect 6787 -581 6887 -547
<< locali >>
rect -6903 547 -6887 581
rect -6787 547 -6771 581
rect -6645 547 -6629 581
rect -6529 547 -6513 581
rect -6387 547 -6371 581
rect -6271 547 -6255 581
rect -6129 547 -6113 581
rect -6013 547 -5997 581
rect -5871 547 -5855 581
rect -5755 547 -5739 581
rect -5613 547 -5597 581
rect -5497 547 -5481 581
rect -5355 547 -5339 581
rect -5239 547 -5223 581
rect -5097 547 -5081 581
rect -4981 547 -4965 581
rect -4839 547 -4823 581
rect -4723 547 -4707 581
rect -4581 547 -4565 581
rect -4465 547 -4449 581
rect -4323 547 -4307 581
rect -4207 547 -4191 581
rect -4065 547 -4049 581
rect -3949 547 -3933 581
rect -3807 547 -3791 581
rect -3691 547 -3675 581
rect -3549 547 -3533 581
rect -3433 547 -3417 581
rect -3291 547 -3275 581
rect -3175 547 -3159 581
rect -3033 547 -3017 581
rect -2917 547 -2901 581
rect -2775 547 -2759 581
rect -2659 547 -2643 581
rect -2517 547 -2501 581
rect -2401 547 -2385 581
rect -2259 547 -2243 581
rect -2143 547 -2127 581
rect -2001 547 -1985 581
rect -1885 547 -1869 581
rect -1743 547 -1727 581
rect -1627 547 -1611 581
rect -1485 547 -1469 581
rect -1369 547 -1353 581
rect -1227 547 -1211 581
rect -1111 547 -1095 581
rect -969 547 -953 581
rect -853 547 -837 581
rect -711 547 -695 581
rect -595 547 -579 581
rect -453 547 -437 581
rect -337 547 -321 581
rect -195 547 -179 581
rect -79 547 -63 581
rect 63 547 79 581
rect 179 547 195 581
rect 321 547 337 581
rect 437 547 453 581
rect 579 547 595 581
rect 695 547 711 581
rect 837 547 853 581
rect 953 547 969 581
rect 1095 547 1111 581
rect 1211 547 1227 581
rect 1353 547 1369 581
rect 1469 547 1485 581
rect 1611 547 1627 581
rect 1727 547 1743 581
rect 1869 547 1885 581
rect 1985 547 2001 581
rect 2127 547 2143 581
rect 2243 547 2259 581
rect 2385 547 2401 581
rect 2501 547 2517 581
rect 2643 547 2659 581
rect 2759 547 2775 581
rect 2901 547 2917 581
rect 3017 547 3033 581
rect 3159 547 3175 581
rect 3275 547 3291 581
rect 3417 547 3433 581
rect 3533 547 3549 581
rect 3675 547 3691 581
rect 3791 547 3807 581
rect 3933 547 3949 581
rect 4049 547 4065 581
rect 4191 547 4207 581
rect 4307 547 4323 581
rect 4449 547 4465 581
rect 4565 547 4581 581
rect 4707 547 4723 581
rect 4823 547 4839 581
rect 4965 547 4981 581
rect 5081 547 5097 581
rect 5223 547 5239 581
rect 5339 547 5355 581
rect 5481 547 5497 581
rect 5597 547 5613 581
rect 5739 547 5755 581
rect 5855 547 5871 581
rect 5997 547 6013 581
rect 6113 547 6129 581
rect 6255 547 6271 581
rect 6371 547 6387 581
rect 6513 547 6529 581
rect 6629 547 6645 581
rect 6771 547 6787 581
rect 6887 547 6903 581
rect -6983 488 -6949 504
rect -6983 -504 -6949 -488
rect -6725 488 -6691 504
rect -6725 -504 -6691 -488
rect -6467 488 -6433 504
rect -6467 -504 -6433 -488
rect -6209 488 -6175 504
rect -6209 -504 -6175 -488
rect -5951 488 -5917 504
rect -5951 -504 -5917 -488
rect -5693 488 -5659 504
rect -5693 -504 -5659 -488
rect -5435 488 -5401 504
rect -5435 -504 -5401 -488
rect -5177 488 -5143 504
rect -5177 -504 -5143 -488
rect -4919 488 -4885 504
rect -4919 -504 -4885 -488
rect -4661 488 -4627 504
rect -4661 -504 -4627 -488
rect -4403 488 -4369 504
rect -4403 -504 -4369 -488
rect -4145 488 -4111 504
rect -4145 -504 -4111 -488
rect -3887 488 -3853 504
rect -3887 -504 -3853 -488
rect -3629 488 -3595 504
rect -3629 -504 -3595 -488
rect -3371 488 -3337 504
rect -3371 -504 -3337 -488
rect -3113 488 -3079 504
rect -3113 -504 -3079 -488
rect -2855 488 -2821 504
rect -2855 -504 -2821 -488
rect -2597 488 -2563 504
rect -2597 -504 -2563 -488
rect -2339 488 -2305 504
rect -2339 -504 -2305 -488
rect -2081 488 -2047 504
rect -2081 -504 -2047 -488
rect -1823 488 -1789 504
rect -1823 -504 -1789 -488
rect -1565 488 -1531 504
rect -1565 -504 -1531 -488
rect -1307 488 -1273 504
rect -1307 -504 -1273 -488
rect -1049 488 -1015 504
rect -1049 -504 -1015 -488
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -504 1049 -488
rect 1273 488 1307 504
rect 1273 -504 1307 -488
rect 1531 488 1565 504
rect 1531 -504 1565 -488
rect 1789 488 1823 504
rect 1789 -504 1823 -488
rect 2047 488 2081 504
rect 2047 -504 2081 -488
rect 2305 488 2339 504
rect 2305 -504 2339 -488
rect 2563 488 2597 504
rect 2563 -504 2597 -488
rect 2821 488 2855 504
rect 2821 -504 2855 -488
rect 3079 488 3113 504
rect 3079 -504 3113 -488
rect 3337 488 3371 504
rect 3337 -504 3371 -488
rect 3595 488 3629 504
rect 3595 -504 3629 -488
rect 3853 488 3887 504
rect 3853 -504 3887 -488
rect 4111 488 4145 504
rect 4111 -504 4145 -488
rect 4369 488 4403 504
rect 4369 -504 4403 -488
rect 4627 488 4661 504
rect 4627 -504 4661 -488
rect 4885 488 4919 504
rect 4885 -504 4919 -488
rect 5143 488 5177 504
rect 5143 -504 5177 -488
rect 5401 488 5435 504
rect 5401 -504 5435 -488
rect 5659 488 5693 504
rect 5659 -504 5693 -488
rect 5917 488 5951 504
rect 5917 -504 5951 -488
rect 6175 488 6209 504
rect 6175 -504 6209 -488
rect 6433 488 6467 504
rect 6433 -504 6467 -488
rect 6691 488 6725 504
rect 6691 -504 6725 -488
rect 6949 488 6983 504
rect 6949 -504 6983 -488
rect -6903 -581 -6887 -547
rect -6787 -581 -6771 -547
rect -6645 -581 -6629 -547
rect -6529 -581 -6513 -547
rect -6387 -581 -6371 -547
rect -6271 -581 -6255 -547
rect -6129 -581 -6113 -547
rect -6013 -581 -5997 -547
rect -5871 -581 -5855 -547
rect -5755 -581 -5739 -547
rect -5613 -581 -5597 -547
rect -5497 -581 -5481 -547
rect -5355 -581 -5339 -547
rect -5239 -581 -5223 -547
rect -5097 -581 -5081 -547
rect -4981 -581 -4965 -547
rect -4839 -581 -4823 -547
rect -4723 -581 -4707 -547
rect -4581 -581 -4565 -547
rect -4465 -581 -4449 -547
rect -4323 -581 -4307 -547
rect -4207 -581 -4191 -547
rect -4065 -581 -4049 -547
rect -3949 -581 -3933 -547
rect -3807 -581 -3791 -547
rect -3691 -581 -3675 -547
rect -3549 -581 -3533 -547
rect -3433 -581 -3417 -547
rect -3291 -581 -3275 -547
rect -3175 -581 -3159 -547
rect -3033 -581 -3017 -547
rect -2917 -581 -2901 -547
rect -2775 -581 -2759 -547
rect -2659 -581 -2643 -547
rect -2517 -581 -2501 -547
rect -2401 -581 -2385 -547
rect -2259 -581 -2243 -547
rect -2143 -581 -2127 -547
rect -2001 -581 -1985 -547
rect -1885 -581 -1869 -547
rect -1743 -581 -1727 -547
rect -1627 -581 -1611 -547
rect -1485 -581 -1469 -547
rect -1369 -581 -1353 -547
rect -1227 -581 -1211 -547
rect -1111 -581 -1095 -547
rect -969 -581 -953 -547
rect -853 -581 -837 -547
rect -711 -581 -695 -547
rect -595 -581 -579 -547
rect -453 -581 -437 -547
rect -337 -581 -321 -547
rect -195 -581 -179 -547
rect -79 -581 -63 -547
rect 63 -581 79 -547
rect 179 -581 195 -547
rect 321 -581 337 -547
rect 437 -581 453 -547
rect 579 -581 595 -547
rect 695 -581 711 -547
rect 837 -581 853 -547
rect 953 -581 969 -547
rect 1095 -581 1111 -547
rect 1211 -581 1227 -547
rect 1353 -581 1369 -547
rect 1469 -581 1485 -547
rect 1611 -581 1627 -547
rect 1727 -581 1743 -547
rect 1869 -581 1885 -547
rect 1985 -581 2001 -547
rect 2127 -581 2143 -547
rect 2243 -581 2259 -547
rect 2385 -581 2401 -547
rect 2501 -581 2517 -547
rect 2643 -581 2659 -547
rect 2759 -581 2775 -547
rect 2901 -581 2917 -547
rect 3017 -581 3033 -547
rect 3159 -581 3175 -547
rect 3275 -581 3291 -547
rect 3417 -581 3433 -547
rect 3533 -581 3549 -547
rect 3675 -581 3691 -547
rect 3791 -581 3807 -547
rect 3933 -581 3949 -547
rect 4049 -581 4065 -547
rect 4191 -581 4207 -547
rect 4307 -581 4323 -547
rect 4449 -581 4465 -547
rect 4565 -581 4581 -547
rect 4707 -581 4723 -547
rect 4823 -581 4839 -547
rect 4965 -581 4981 -547
rect 5081 -581 5097 -547
rect 5223 -581 5239 -547
rect 5339 -581 5355 -547
rect 5481 -581 5497 -547
rect 5597 -581 5613 -547
rect 5739 -581 5755 -547
rect 5855 -581 5871 -547
rect 5997 -581 6013 -547
rect 6113 -581 6129 -547
rect 6255 -581 6271 -547
rect 6371 -581 6387 -547
rect 6513 -581 6529 -547
rect 6629 -581 6645 -547
rect 6771 -581 6787 -547
rect 6887 -581 6903 -547
<< viali >>
rect -6871 547 -6803 581
rect -6613 547 -6545 581
rect -6355 547 -6287 581
rect -6097 547 -6029 581
rect -5839 547 -5771 581
rect -5581 547 -5513 581
rect -5323 547 -5255 581
rect -5065 547 -4997 581
rect -4807 547 -4739 581
rect -4549 547 -4481 581
rect -4291 547 -4223 581
rect -4033 547 -3965 581
rect -3775 547 -3707 581
rect -3517 547 -3449 581
rect -3259 547 -3191 581
rect -3001 547 -2933 581
rect -2743 547 -2675 581
rect -2485 547 -2417 581
rect -2227 547 -2159 581
rect -1969 547 -1901 581
rect -1711 547 -1643 581
rect -1453 547 -1385 581
rect -1195 547 -1127 581
rect -937 547 -869 581
rect -679 547 -611 581
rect -421 547 -353 581
rect -163 547 -95 581
rect 95 547 163 581
rect 353 547 421 581
rect 611 547 679 581
rect 869 547 937 581
rect 1127 547 1195 581
rect 1385 547 1453 581
rect 1643 547 1711 581
rect 1901 547 1969 581
rect 2159 547 2227 581
rect 2417 547 2485 581
rect 2675 547 2743 581
rect 2933 547 3001 581
rect 3191 547 3259 581
rect 3449 547 3517 581
rect 3707 547 3775 581
rect 3965 547 4033 581
rect 4223 547 4291 581
rect 4481 547 4549 581
rect 4739 547 4807 581
rect 4997 547 5065 581
rect 5255 547 5323 581
rect 5513 547 5581 581
rect 5771 547 5839 581
rect 6029 547 6097 581
rect 6287 547 6355 581
rect 6545 547 6613 581
rect 6803 547 6871 581
rect -6983 -488 -6949 488
rect -6725 -488 -6691 488
rect -6467 -488 -6433 488
rect -6209 -488 -6175 488
rect -5951 -488 -5917 488
rect -5693 -488 -5659 488
rect -5435 -488 -5401 488
rect -5177 -488 -5143 488
rect -4919 -488 -4885 488
rect -4661 -488 -4627 488
rect -4403 -488 -4369 488
rect -4145 -488 -4111 488
rect -3887 -488 -3853 488
rect -3629 -488 -3595 488
rect -3371 -488 -3337 488
rect -3113 -488 -3079 488
rect -2855 -488 -2821 488
rect -2597 -488 -2563 488
rect -2339 -488 -2305 488
rect -2081 -488 -2047 488
rect -1823 -488 -1789 488
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect 1789 -488 1823 488
rect 2047 -488 2081 488
rect 2305 -488 2339 488
rect 2563 -488 2597 488
rect 2821 -488 2855 488
rect 3079 -488 3113 488
rect 3337 -488 3371 488
rect 3595 -488 3629 488
rect 3853 -488 3887 488
rect 4111 -488 4145 488
rect 4369 -488 4403 488
rect 4627 -488 4661 488
rect 4885 -488 4919 488
rect 5143 -488 5177 488
rect 5401 -488 5435 488
rect 5659 -488 5693 488
rect 5917 -488 5951 488
rect 6175 -488 6209 488
rect 6433 -488 6467 488
rect 6691 -488 6725 488
rect 6949 -488 6983 488
rect -6871 -581 -6803 -547
rect -6613 -581 -6545 -547
rect -6355 -581 -6287 -547
rect -6097 -581 -6029 -547
rect -5839 -581 -5771 -547
rect -5581 -581 -5513 -547
rect -5323 -581 -5255 -547
rect -5065 -581 -4997 -547
rect -4807 -581 -4739 -547
rect -4549 -581 -4481 -547
rect -4291 -581 -4223 -547
rect -4033 -581 -3965 -547
rect -3775 -581 -3707 -547
rect -3517 -581 -3449 -547
rect -3259 -581 -3191 -547
rect -3001 -581 -2933 -547
rect -2743 -581 -2675 -547
rect -2485 -581 -2417 -547
rect -2227 -581 -2159 -547
rect -1969 -581 -1901 -547
rect -1711 -581 -1643 -547
rect -1453 -581 -1385 -547
rect -1195 -581 -1127 -547
rect -937 -581 -869 -547
rect -679 -581 -611 -547
rect -421 -581 -353 -547
rect -163 -581 -95 -547
rect 95 -581 163 -547
rect 353 -581 421 -547
rect 611 -581 679 -547
rect 869 -581 937 -547
rect 1127 -581 1195 -547
rect 1385 -581 1453 -547
rect 1643 -581 1711 -547
rect 1901 -581 1969 -547
rect 2159 -581 2227 -547
rect 2417 -581 2485 -547
rect 2675 -581 2743 -547
rect 2933 -581 3001 -547
rect 3191 -581 3259 -547
rect 3449 -581 3517 -547
rect 3707 -581 3775 -547
rect 3965 -581 4033 -547
rect 4223 -581 4291 -547
rect 4481 -581 4549 -547
rect 4739 -581 4807 -547
rect 4997 -581 5065 -547
rect 5255 -581 5323 -547
rect 5513 -581 5581 -547
rect 5771 -581 5839 -547
rect 6029 -581 6097 -547
rect 6287 -581 6355 -547
rect 6545 -581 6613 -547
rect 6803 -581 6871 -547
<< metal1 >>
rect -6883 581 -6791 587
rect -6883 547 -6871 581
rect -6803 547 -6791 581
rect -6883 541 -6791 547
rect -6625 581 -6533 587
rect -6625 547 -6613 581
rect -6545 547 -6533 581
rect -6625 541 -6533 547
rect -6367 581 -6275 587
rect -6367 547 -6355 581
rect -6287 547 -6275 581
rect -6367 541 -6275 547
rect -6109 581 -6017 587
rect -6109 547 -6097 581
rect -6029 547 -6017 581
rect -6109 541 -6017 547
rect -5851 581 -5759 587
rect -5851 547 -5839 581
rect -5771 547 -5759 581
rect -5851 541 -5759 547
rect -5593 581 -5501 587
rect -5593 547 -5581 581
rect -5513 547 -5501 581
rect -5593 541 -5501 547
rect -5335 581 -5243 587
rect -5335 547 -5323 581
rect -5255 547 -5243 581
rect -5335 541 -5243 547
rect -5077 581 -4985 587
rect -5077 547 -5065 581
rect -4997 547 -4985 581
rect -5077 541 -4985 547
rect -4819 581 -4727 587
rect -4819 547 -4807 581
rect -4739 547 -4727 581
rect -4819 541 -4727 547
rect -4561 581 -4469 587
rect -4561 547 -4549 581
rect -4481 547 -4469 581
rect -4561 541 -4469 547
rect -4303 581 -4211 587
rect -4303 547 -4291 581
rect -4223 547 -4211 581
rect -4303 541 -4211 547
rect -4045 581 -3953 587
rect -4045 547 -4033 581
rect -3965 547 -3953 581
rect -4045 541 -3953 547
rect -3787 581 -3695 587
rect -3787 547 -3775 581
rect -3707 547 -3695 581
rect -3787 541 -3695 547
rect -3529 581 -3437 587
rect -3529 547 -3517 581
rect -3449 547 -3437 581
rect -3529 541 -3437 547
rect -3271 581 -3179 587
rect -3271 547 -3259 581
rect -3191 547 -3179 581
rect -3271 541 -3179 547
rect -3013 581 -2921 587
rect -3013 547 -3001 581
rect -2933 547 -2921 581
rect -3013 541 -2921 547
rect -2755 581 -2663 587
rect -2755 547 -2743 581
rect -2675 547 -2663 581
rect -2755 541 -2663 547
rect -2497 581 -2405 587
rect -2497 547 -2485 581
rect -2417 547 -2405 581
rect -2497 541 -2405 547
rect -2239 581 -2147 587
rect -2239 547 -2227 581
rect -2159 547 -2147 581
rect -2239 541 -2147 547
rect -1981 581 -1889 587
rect -1981 547 -1969 581
rect -1901 547 -1889 581
rect -1981 541 -1889 547
rect -1723 581 -1631 587
rect -1723 547 -1711 581
rect -1643 547 -1631 581
rect -1723 541 -1631 547
rect -1465 581 -1373 587
rect -1465 547 -1453 581
rect -1385 547 -1373 581
rect -1465 541 -1373 547
rect -1207 581 -1115 587
rect -1207 547 -1195 581
rect -1127 547 -1115 581
rect -1207 541 -1115 547
rect -949 581 -857 587
rect -949 547 -937 581
rect -869 547 -857 581
rect -949 541 -857 547
rect -691 581 -599 587
rect -691 547 -679 581
rect -611 547 -599 581
rect -691 541 -599 547
rect -433 581 -341 587
rect -433 547 -421 581
rect -353 547 -341 581
rect -433 541 -341 547
rect -175 581 -83 587
rect -175 547 -163 581
rect -95 547 -83 581
rect -175 541 -83 547
rect 83 581 175 587
rect 83 547 95 581
rect 163 547 175 581
rect 83 541 175 547
rect 341 581 433 587
rect 341 547 353 581
rect 421 547 433 581
rect 341 541 433 547
rect 599 581 691 587
rect 599 547 611 581
rect 679 547 691 581
rect 599 541 691 547
rect 857 581 949 587
rect 857 547 869 581
rect 937 547 949 581
rect 857 541 949 547
rect 1115 581 1207 587
rect 1115 547 1127 581
rect 1195 547 1207 581
rect 1115 541 1207 547
rect 1373 581 1465 587
rect 1373 547 1385 581
rect 1453 547 1465 581
rect 1373 541 1465 547
rect 1631 581 1723 587
rect 1631 547 1643 581
rect 1711 547 1723 581
rect 1631 541 1723 547
rect 1889 581 1981 587
rect 1889 547 1901 581
rect 1969 547 1981 581
rect 1889 541 1981 547
rect 2147 581 2239 587
rect 2147 547 2159 581
rect 2227 547 2239 581
rect 2147 541 2239 547
rect 2405 581 2497 587
rect 2405 547 2417 581
rect 2485 547 2497 581
rect 2405 541 2497 547
rect 2663 581 2755 587
rect 2663 547 2675 581
rect 2743 547 2755 581
rect 2663 541 2755 547
rect 2921 581 3013 587
rect 2921 547 2933 581
rect 3001 547 3013 581
rect 2921 541 3013 547
rect 3179 581 3271 587
rect 3179 547 3191 581
rect 3259 547 3271 581
rect 3179 541 3271 547
rect 3437 581 3529 587
rect 3437 547 3449 581
rect 3517 547 3529 581
rect 3437 541 3529 547
rect 3695 581 3787 587
rect 3695 547 3707 581
rect 3775 547 3787 581
rect 3695 541 3787 547
rect 3953 581 4045 587
rect 3953 547 3965 581
rect 4033 547 4045 581
rect 3953 541 4045 547
rect 4211 581 4303 587
rect 4211 547 4223 581
rect 4291 547 4303 581
rect 4211 541 4303 547
rect 4469 581 4561 587
rect 4469 547 4481 581
rect 4549 547 4561 581
rect 4469 541 4561 547
rect 4727 581 4819 587
rect 4727 547 4739 581
rect 4807 547 4819 581
rect 4727 541 4819 547
rect 4985 581 5077 587
rect 4985 547 4997 581
rect 5065 547 5077 581
rect 4985 541 5077 547
rect 5243 581 5335 587
rect 5243 547 5255 581
rect 5323 547 5335 581
rect 5243 541 5335 547
rect 5501 581 5593 587
rect 5501 547 5513 581
rect 5581 547 5593 581
rect 5501 541 5593 547
rect 5759 581 5851 587
rect 5759 547 5771 581
rect 5839 547 5851 581
rect 5759 541 5851 547
rect 6017 581 6109 587
rect 6017 547 6029 581
rect 6097 547 6109 581
rect 6017 541 6109 547
rect 6275 581 6367 587
rect 6275 547 6287 581
rect 6355 547 6367 581
rect 6275 541 6367 547
rect 6533 581 6625 587
rect 6533 547 6545 581
rect 6613 547 6625 581
rect 6533 541 6625 547
rect 6791 581 6883 587
rect 6791 547 6803 581
rect 6871 547 6883 581
rect 6791 541 6883 547
rect -6989 488 -6943 500
rect -6989 -488 -6983 488
rect -6949 -488 -6943 488
rect -6989 -500 -6943 -488
rect -6731 488 -6685 500
rect -6731 -488 -6725 488
rect -6691 -488 -6685 488
rect -6731 -500 -6685 -488
rect -6473 488 -6427 500
rect -6473 -488 -6467 488
rect -6433 -488 -6427 488
rect -6473 -500 -6427 -488
rect -6215 488 -6169 500
rect -6215 -488 -6209 488
rect -6175 -488 -6169 488
rect -6215 -500 -6169 -488
rect -5957 488 -5911 500
rect -5957 -488 -5951 488
rect -5917 -488 -5911 488
rect -5957 -500 -5911 -488
rect -5699 488 -5653 500
rect -5699 -488 -5693 488
rect -5659 -488 -5653 488
rect -5699 -500 -5653 -488
rect -5441 488 -5395 500
rect -5441 -488 -5435 488
rect -5401 -488 -5395 488
rect -5441 -500 -5395 -488
rect -5183 488 -5137 500
rect -5183 -488 -5177 488
rect -5143 -488 -5137 488
rect -5183 -500 -5137 -488
rect -4925 488 -4879 500
rect -4925 -488 -4919 488
rect -4885 -488 -4879 488
rect -4925 -500 -4879 -488
rect -4667 488 -4621 500
rect -4667 -488 -4661 488
rect -4627 -488 -4621 488
rect -4667 -500 -4621 -488
rect -4409 488 -4363 500
rect -4409 -488 -4403 488
rect -4369 -488 -4363 488
rect -4409 -500 -4363 -488
rect -4151 488 -4105 500
rect -4151 -488 -4145 488
rect -4111 -488 -4105 488
rect -4151 -500 -4105 -488
rect -3893 488 -3847 500
rect -3893 -488 -3887 488
rect -3853 -488 -3847 488
rect -3893 -500 -3847 -488
rect -3635 488 -3589 500
rect -3635 -488 -3629 488
rect -3595 -488 -3589 488
rect -3635 -500 -3589 -488
rect -3377 488 -3331 500
rect -3377 -488 -3371 488
rect -3337 -488 -3331 488
rect -3377 -500 -3331 -488
rect -3119 488 -3073 500
rect -3119 -488 -3113 488
rect -3079 -488 -3073 488
rect -3119 -500 -3073 -488
rect -2861 488 -2815 500
rect -2861 -488 -2855 488
rect -2821 -488 -2815 488
rect -2861 -500 -2815 -488
rect -2603 488 -2557 500
rect -2603 -488 -2597 488
rect -2563 -488 -2557 488
rect -2603 -500 -2557 -488
rect -2345 488 -2299 500
rect -2345 -488 -2339 488
rect -2305 -488 -2299 488
rect -2345 -500 -2299 -488
rect -2087 488 -2041 500
rect -2087 -488 -2081 488
rect -2047 -488 -2041 488
rect -2087 -500 -2041 -488
rect -1829 488 -1783 500
rect -1829 -488 -1823 488
rect -1789 -488 -1783 488
rect -1829 -500 -1783 -488
rect -1571 488 -1525 500
rect -1571 -488 -1565 488
rect -1531 -488 -1525 488
rect -1571 -500 -1525 -488
rect -1313 488 -1267 500
rect -1313 -488 -1307 488
rect -1273 -488 -1267 488
rect -1313 -500 -1267 -488
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect 1267 488 1313 500
rect 1267 -488 1273 488
rect 1307 -488 1313 488
rect 1267 -500 1313 -488
rect 1525 488 1571 500
rect 1525 -488 1531 488
rect 1565 -488 1571 488
rect 1525 -500 1571 -488
rect 1783 488 1829 500
rect 1783 -488 1789 488
rect 1823 -488 1829 488
rect 1783 -500 1829 -488
rect 2041 488 2087 500
rect 2041 -488 2047 488
rect 2081 -488 2087 488
rect 2041 -500 2087 -488
rect 2299 488 2345 500
rect 2299 -488 2305 488
rect 2339 -488 2345 488
rect 2299 -500 2345 -488
rect 2557 488 2603 500
rect 2557 -488 2563 488
rect 2597 -488 2603 488
rect 2557 -500 2603 -488
rect 2815 488 2861 500
rect 2815 -488 2821 488
rect 2855 -488 2861 488
rect 2815 -500 2861 -488
rect 3073 488 3119 500
rect 3073 -488 3079 488
rect 3113 -488 3119 488
rect 3073 -500 3119 -488
rect 3331 488 3377 500
rect 3331 -488 3337 488
rect 3371 -488 3377 488
rect 3331 -500 3377 -488
rect 3589 488 3635 500
rect 3589 -488 3595 488
rect 3629 -488 3635 488
rect 3589 -500 3635 -488
rect 3847 488 3893 500
rect 3847 -488 3853 488
rect 3887 -488 3893 488
rect 3847 -500 3893 -488
rect 4105 488 4151 500
rect 4105 -488 4111 488
rect 4145 -488 4151 488
rect 4105 -500 4151 -488
rect 4363 488 4409 500
rect 4363 -488 4369 488
rect 4403 -488 4409 488
rect 4363 -500 4409 -488
rect 4621 488 4667 500
rect 4621 -488 4627 488
rect 4661 -488 4667 488
rect 4621 -500 4667 -488
rect 4879 488 4925 500
rect 4879 -488 4885 488
rect 4919 -488 4925 488
rect 4879 -500 4925 -488
rect 5137 488 5183 500
rect 5137 -488 5143 488
rect 5177 -488 5183 488
rect 5137 -500 5183 -488
rect 5395 488 5441 500
rect 5395 -488 5401 488
rect 5435 -488 5441 488
rect 5395 -500 5441 -488
rect 5653 488 5699 500
rect 5653 -488 5659 488
rect 5693 -488 5699 488
rect 5653 -500 5699 -488
rect 5911 488 5957 500
rect 5911 -488 5917 488
rect 5951 -488 5957 488
rect 5911 -500 5957 -488
rect 6169 488 6215 500
rect 6169 -488 6175 488
rect 6209 -488 6215 488
rect 6169 -500 6215 -488
rect 6427 488 6473 500
rect 6427 -488 6433 488
rect 6467 -488 6473 488
rect 6427 -500 6473 -488
rect 6685 488 6731 500
rect 6685 -488 6691 488
rect 6725 -488 6731 488
rect 6685 -500 6731 -488
rect 6943 488 6989 500
rect 6943 -488 6949 488
rect 6983 -488 6989 488
rect 6943 -500 6989 -488
rect -6883 -547 -6791 -541
rect -6883 -581 -6871 -547
rect -6803 -581 -6791 -547
rect -6883 -587 -6791 -581
rect -6625 -547 -6533 -541
rect -6625 -581 -6613 -547
rect -6545 -581 -6533 -547
rect -6625 -587 -6533 -581
rect -6367 -547 -6275 -541
rect -6367 -581 -6355 -547
rect -6287 -581 -6275 -547
rect -6367 -587 -6275 -581
rect -6109 -547 -6017 -541
rect -6109 -581 -6097 -547
rect -6029 -581 -6017 -547
rect -6109 -587 -6017 -581
rect -5851 -547 -5759 -541
rect -5851 -581 -5839 -547
rect -5771 -581 -5759 -547
rect -5851 -587 -5759 -581
rect -5593 -547 -5501 -541
rect -5593 -581 -5581 -547
rect -5513 -581 -5501 -547
rect -5593 -587 -5501 -581
rect -5335 -547 -5243 -541
rect -5335 -581 -5323 -547
rect -5255 -581 -5243 -547
rect -5335 -587 -5243 -581
rect -5077 -547 -4985 -541
rect -5077 -581 -5065 -547
rect -4997 -581 -4985 -547
rect -5077 -587 -4985 -581
rect -4819 -547 -4727 -541
rect -4819 -581 -4807 -547
rect -4739 -581 -4727 -547
rect -4819 -587 -4727 -581
rect -4561 -547 -4469 -541
rect -4561 -581 -4549 -547
rect -4481 -581 -4469 -547
rect -4561 -587 -4469 -581
rect -4303 -547 -4211 -541
rect -4303 -581 -4291 -547
rect -4223 -581 -4211 -547
rect -4303 -587 -4211 -581
rect -4045 -547 -3953 -541
rect -4045 -581 -4033 -547
rect -3965 -581 -3953 -547
rect -4045 -587 -3953 -581
rect -3787 -547 -3695 -541
rect -3787 -581 -3775 -547
rect -3707 -581 -3695 -547
rect -3787 -587 -3695 -581
rect -3529 -547 -3437 -541
rect -3529 -581 -3517 -547
rect -3449 -581 -3437 -547
rect -3529 -587 -3437 -581
rect -3271 -547 -3179 -541
rect -3271 -581 -3259 -547
rect -3191 -581 -3179 -547
rect -3271 -587 -3179 -581
rect -3013 -547 -2921 -541
rect -3013 -581 -3001 -547
rect -2933 -581 -2921 -547
rect -3013 -587 -2921 -581
rect -2755 -547 -2663 -541
rect -2755 -581 -2743 -547
rect -2675 -581 -2663 -547
rect -2755 -587 -2663 -581
rect -2497 -547 -2405 -541
rect -2497 -581 -2485 -547
rect -2417 -581 -2405 -547
rect -2497 -587 -2405 -581
rect -2239 -547 -2147 -541
rect -2239 -581 -2227 -547
rect -2159 -581 -2147 -547
rect -2239 -587 -2147 -581
rect -1981 -547 -1889 -541
rect -1981 -581 -1969 -547
rect -1901 -581 -1889 -547
rect -1981 -587 -1889 -581
rect -1723 -547 -1631 -541
rect -1723 -581 -1711 -547
rect -1643 -581 -1631 -547
rect -1723 -587 -1631 -581
rect -1465 -547 -1373 -541
rect -1465 -581 -1453 -547
rect -1385 -581 -1373 -547
rect -1465 -587 -1373 -581
rect -1207 -547 -1115 -541
rect -1207 -581 -1195 -547
rect -1127 -581 -1115 -547
rect -1207 -587 -1115 -581
rect -949 -547 -857 -541
rect -949 -581 -937 -547
rect -869 -581 -857 -547
rect -949 -587 -857 -581
rect -691 -547 -599 -541
rect -691 -581 -679 -547
rect -611 -581 -599 -547
rect -691 -587 -599 -581
rect -433 -547 -341 -541
rect -433 -581 -421 -547
rect -353 -581 -341 -547
rect -433 -587 -341 -581
rect -175 -547 -83 -541
rect -175 -581 -163 -547
rect -95 -581 -83 -547
rect -175 -587 -83 -581
rect 83 -547 175 -541
rect 83 -581 95 -547
rect 163 -581 175 -547
rect 83 -587 175 -581
rect 341 -547 433 -541
rect 341 -581 353 -547
rect 421 -581 433 -547
rect 341 -587 433 -581
rect 599 -547 691 -541
rect 599 -581 611 -547
rect 679 -581 691 -547
rect 599 -587 691 -581
rect 857 -547 949 -541
rect 857 -581 869 -547
rect 937 -581 949 -547
rect 857 -587 949 -581
rect 1115 -547 1207 -541
rect 1115 -581 1127 -547
rect 1195 -581 1207 -547
rect 1115 -587 1207 -581
rect 1373 -547 1465 -541
rect 1373 -581 1385 -547
rect 1453 -581 1465 -547
rect 1373 -587 1465 -581
rect 1631 -547 1723 -541
rect 1631 -581 1643 -547
rect 1711 -581 1723 -547
rect 1631 -587 1723 -581
rect 1889 -547 1981 -541
rect 1889 -581 1901 -547
rect 1969 -581 1981 -547
rect 1889 -587 1981 -581
rect 2147 -547 2239 -541
rect 2147 -581 2159 -547
rect 2227 -581 2239 -547
rect 2147 -587 2239 -581
rect 2405 -547 2497 -541
rect 2405 -581 2417 -547
rect 2485 -581 2497 -547
rect 2405 -587 2497 -581
rect 2663 -547 2755 -541
rect 2663 -581 2675 -547
rect 2743 -581 2755 -547
rect 2663 -587 2755 -581
rect 2921 -547 3013 -541
rect 2921 -581 2933 -547
rect 3001 -581 3013 -547
rect 2921 -587 3013 -581
rect 3179 -547 3271 -541
rect 3179 -581 3191 -547
rect 3259 -581 3271 -547
rect 3179 -587 3271 -581
rect 3437 -547 3529 -541
rect 3437 -581 3449 -547
rect 3517 -581 3529 -547
rect 3437 -587 3529 -581
rect 3695 -547 3787 -541
rect 3695 -581 3707 -547
rect 3775 -581 3787 -547
rect 3695 -587 3787 -581
rect 3953 -547 4045 -541
rect 3953 -581 3965 -547
rect 4033 -581 4045 -547
rect 3953 -587 4045 -581
rect 4211 -547 4303 -541
rect 4211 -581 4223 -547
rect 4291 -581 4303 -547
rect 4211 -587 4303 -581
rect 4469 -547 4561 -541
rect 4469 -581 4481 -547
rect 4549 -581 4561 -547
rect 4469 -587 4561 -581
rect 4727 -547 4819 -541
rect 4727 -581 4739 -547
rect 4807 -581 4819 -547
rect 4727 -587 4819 -581
rect 4985 -547 5077 -541
rect 4985 -581 4997 -547
rect 5065 -581 5077 -547
rect 4985 -587 5077 -581
rect 5243 -547 5335 -541
rect 5243 -581 5255 -547
rect 5323 -581 5335 -547
rect 5243 -587 5335 -581
rect 5501 -547 5593 -541
rect 5501 -581 5513 -547
rect 5581 -581 5593 -547
rect 5501 -587 5593 -581
rect 5759 -547 5851 -541
rect 5759 -581 5771 -547
rect 5839 -581 5851 -547
rect 5759 -587 5851 -581
rect 6017 -547 6109 -541
rect 6017 -581 6029 -547
rect 6097 -581 6109 -547
rect 6017 -587 6109 -581
rect 6275 -547 6367 -541
rect 6275 -581 6287 -547
rect 6355 -581 6367 -547
rect 6275 -587 6367 -581
rect 6533 -547 6625 -541
rect 6533 -581 6545 -547
rect 6613 -581 6625 -547
rect 6533 -587 6625 -581
rect 6791 -547 6883 -541
rect 6791 -581 6803 -547
rect 6871 -581 6883 -547
rect 6791 -587 6883 -581
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string parameters w 5 l 1 m 1 nf 54 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
