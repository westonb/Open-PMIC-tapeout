magic
tech sky130A
magscale 1 2
timestamp 1624002729
<< nwell >>
rect -3000 40 3000 4500
<< pwell >>
rect -3000 -4500 3000 -40
<< mvnmos >>
rect -1677 -1700 -1477 -700
rect -1419 -1700 -1319 -700
rect -1261 -1700 -1061 -700
rect -1003 -1700 -803 -700
rect -745 -1700 -545 -700
rect -487 -1700 -287 -700
rect -229 -1700 -29 -700
rect 29 -1700 229 -700
rect 287 -1700 487 -700
rect 545 -1700 745 -700
rect 803 -1700 1003 -700
rect 1061 -1700 1261 -700
rect 1319 -1700 1419 -700
rect 1477 -1700 1677 -700
rect -2293 -3500 -2093 -2500
rect -2035 -3500 -1835 -2500
rect -1777 -3500 -1577 -2500
rect -1519 -3500 -1319 -2500
rect -1261 -3500 -1061 -2500
rect -1003 -3500 -803 -2500
rect -745 -3500 -545 -2500
rect -487 -3500 -287 -2500
rect -229 -3500 -29 -2500
rect 29 -3500 229 -2500
rect 287 -3500 487 -2500
rect 545 -3500 745 -2500
rect 803 -3500 1003 -2500
rect 1061 -3500 1261 -2500
rect 1319 -3500 1519 -2500
rect 1577 -3500 1777 -2500
rect 1835 -3500 2035 -2500
rect 2093 -3500 2293 -2500
<< mvpmos >>
rect -2293 2500 -2093 3500
rect -2035 2500 -1835 3500
rect -1777 2500 -1577 3500
rect -1519 2500 -1319 3500
rect -1261 2500 -1061 3500
rect -1003 2500 -803 3500
rect -745 2500 -545 3500
rect -487 2500 -287 3500
rect -229 2500 -29 3500
rect 29 2500 229 3500
rect 287 2500 487 3500
rect 545 2500 745 3500
rect 803 2500 1003 3500
rect 1061 2500 1261 3500
rect 1319 2500 1519 3500
rect 1577 2500 1777 3500
rect 1835 2500 2035 3500
rect 2093 2500 2293 3500
rect -1677 700 -1477 1700
rect -1419 700 -1319 1700
rect -1261 700 -1061 1700
rect -1003 700 -803 1700
rect -745 700 -545 1700
rect -487 700 -287 1700
rect -229 700 -29 1700
rect 29 700 229 1700
rect 287 700 487 1700
rect 545 700 745 1700
rect 803 700 1003 1700
rect 1061 700 1261 1700
rect 1319 700 1419 1700
rect 1477 700 1677 1700
<< mvndiff >>
rect -1735 -712 -1677 -700
rect -1735 -1688 -1723 -712
rect -1689 -1688 -1677 -712
rect -1735 -1700 -1677 -1688
rect -1477 -712 -1419 -700
rect -1477 -1688 -1465 -712
rect -1431 -1688 -1419 -712
rect -1477 -1700 -1419 -1688
rect -1319 -712 -1261 -700
rect -1319 -1688 -1307 -712
rect -1273 -1688 -1261 -712
rect -1319 -1700 -1261 -1688
rect -1061 -712 -1003 -700
rect -1061 -1688 -1049 -712
rect -1015 -1688 -1003 -712
rect -1061 -1700 -1003 -1688
rect -803 -712 -745 -700
rect -803 -1688 -791 -712
rect -757 -1688 -745 -712
rect -803 -1700 -745 -1688
rect -545 -712 -487 -700
rect -545 -1688 -533 -712
rect -499 -1688 -487 -712
rect -545 -1700 -487 -1688
rect -287 -712 -229 -700
rect -287 -1688 -275 -712
rect -241 -1688 -229 -712
rect -287 -1700 -229 -1688
rect -29 -712 29 -700
rect -29 -1688 -17 -712
rect 17 -1688 29 -712
rect -29 -1700 29 -1688
rect 229 -712 287 -700
rect 229 -1688 241 -712
rect 275 -1688 287 -712
rect 229 -1700 287 -1688
rect 487 -712 545 -700
rect 487 -1688 499 -712
rect 533 -1688 545 -712
rect 487 -1700 545 -1688
rect 745 -712 803 -700
rect 745 -1688 757 -712
rect 791 -1688 803 -712
rect 745 -1700 803 -1688
rect 1003 -712 1061 -700
rect 1003 -1688 1015 -712
rect 1049 -1688 1061 -712
rect 1003 -1700 1061 -1688
rect 1261 -712 1319 -700
rect 1261 -1688 1273 -712
rect 1307 -1688 1319 -712
rect 1261 -1700 1319 -1688
rect 1419 -712 1477 -700
rect 1419 -1688 1431 -712
rect 1465 -1688 1477 -712
rect 1419 -1700 1477 -1688
rect 1677 -712 1735 -700
rect 1677 -1688 1689 -712
rect 1723 -1688 1735 -712
rect 1677 -1700 1735 -1688
rect -2351 -2512 -2293 -2500
rect -2351 -3488 -2339 -2512
rect -2305 -3488 -2293 -2512
rect -2351 -3500 -2293 -3488
rect -2093 -2512 -2035 -2500
rect -2093 -3488 -2081 -2512
rect -2047 -3488 -2035 -2512
rect -2093 -3500 -2035 -3488
rect -1835 -2512 -1777 -2500
rect -1835 -3488 -1823 -2512
rect -1789 -3488 -1777 -2512
rect -1835 -3500 -1777 -3488
rect -1577 -2512 -1519 -2500
rect -1577 -3488 -1565 -2512
rect -1531 -3488 -1519 -2512
rect -1577 -3500 -1519 -3488
rect -1319 -2512 -1261 -2500
rect -1319 -3488 -1307 -2512
rect -1273 -3488 -1261 -2512
rect -1319 -3500 -1261 -3488
rect -1061 -2512 -1003 -2500
rect -1061 -3488 -1049 -2512
rect -1015 -3488 -1003 -2512
rect -1061 -3500 -1003 -3488
rect -803 -2512 -745 -2500
rect -803 -3488 -791 -2512
rect -757 -3488 -745 -2512
rect -803 -3500 -745 -3488
rect -545 -2512 -487 -2500
rect -545 -3488 -533 -2512
rect -499 -3488 -487 -2512
rect -545 -3500 -487 -3488
rect -287 -2512 -229 -2500
rect -287 -3488 -275 -2512
rect -241 -3488 -229 -2512
rect -287 -3500 -229 -3488
rect -29 -2512 29 -2500
rect -29 -3488 -17 -2512
rect 17 -3488 29 -2512
rect -29 -3500 29 -3488
rect 229 -2512 287 -2500
rect 229 -3488 241 -2512
rect 275 -3488 287 -2512
rect 229 -3500 287 -3488
rect 487 -2512 545 -2500
rect 487 -3488 499 -2512
rect 533 -3488 545 -2512
rect 487 -3500 545 -3488
rect 745 -2512 803 -2500
rect 745 -3488 757 -2512
rect 791 -3488 803 -2512
rect 745 -3500 803 -3488
rect 1003 -2512 1061 -2500
rect 1003 -3488 1015 -2512
rect 1049 -3488 1061 -2512
rect 1003 -3500 1061 -3488
rect 1261 -2512 1319 -2500
rect 1261 -3488 1273 -2512
rect 1307 -3488 1319 -2512
rect 1261 -3500 1319 -3488
rect 1519 -2512 1577 -2500
rect 1519 -3488 1531 -2512
rect 1565 -3488 1577 -2512
rect 1519 -3500 1577 -3488
rect 1777 -2512 1835 -2500
rect 1777 -3488 1789 -2512
rect 1823 -3488 1835 -2512
rect 1777 -3500 1835 -3488
rect 2035 -2512 2093 -2500
rect 2035 -3488 2047 -2512
rect 2081 -3488 2093 -2512
rect 2035 -3500 2093 -3488
rect 2293 -2512 2351 -2500
rect 2293 -3488 2305 -2512
rect 2339 -3488 2351 -2512
rect 2293 -3500 2351 -3488
<< mvpdiff >>
rect -2351 3488 -2293 3500
rect -2351 2512 -2339 3488
rect -2305 2512 -2293 3488
rect -2351 2500 -2293 2512
rect -2093 3488 -2035 3500
rect -2093 2512 -2081 3488
rect -2047 2512 -2035 3488
rect -2093 2500 -2035 2512
rect -1835 3488 -1777 3500
rect -1835 2512 -1823 3488
rect -1789 2512 -1777 3488
rect -1835 2500 -1777 2512
rect -1577 3488 -1519 3500
rect -1577 2512 -1565 3488
rect -1531 2512 -1519 3488
rect -1577 2500 -1519 2512
rect -1319 3488 -1261 3500
rect -1319 2512 -1307 3488
rect -1273 2512 -1261 3488
rect -1319 2500 -1261 2512
rect -1061 3488 -1003 3500
rect -1061 2512 -1049 3488
rect -1015 2512 -1003 3488
rect -1061 2500 -1003 2512
rect -803 3488 -745 3500
rect -803 2512 -791 3488
rect -757 2512 -745 3488
rect -803 2500 -745 2512
rect -545 3488 -487 3500
rect -545 2512 -533 3488
rect -499 2512 -487 3488
rect -545 2500 -487 2512
rect -287 3488 -229 3500
rect -287 2512 -275 3488
rect -241 2512 -229 3488
rect -287 2500 -229 2512
rect -29 3488 29 3500
rect -29 2512 -17 3488
rect 17 2512 29 3488
rect -29 2500 29 2512
rect 229 3488 287 3500
rect 229 2512 241 3488
rect 275 2512 287 3488
rect 229 2500 287 2512
rect 487 3488 545 3500
rect 487 2512 499 3488
rect 533 2512 545 3488
rect 487 2500 545 2512
rect 745 3488 803 3500
rect 745 2512 757 3488
rect 791 2512 803 3488
rect 745 2500 803 2512
rect 1003 3488 1061 3500
rect 1003 2512 1015 3488
rect 1049 2512 1061 3488
rect 1003 2500 1061 2512
rect 1261 3488 1319 3500
rect 1261 2512 1273 3488
rect 1307 2512 1319 3488
rect 1261 2500 1319 2512
rect 1519 3488 1577 3500
rect 1519 2512 1531 3488
rect 1565 2512 1577 3488
rect 1519 2500 1577 2512
rect 1777 3488 1835 3500
rect 1777 2512 1789 3488
rect 1823 2512 1835 3488
rect 1777 2500 1835 2512
rect 2035 3488 2093 3500
rect 2035 2512 2047 3488
rect 2081 2512 2093 3488
rect 2035 2500 2093 2512
rect 2293 3488 2351 3500
rect 2293 2512 2305 3488
rect 2339 2512 2351 3488
rect 2293 2500 2351 2512
rect -1735 1688 -1677 1700
rect -1735 712 -1723 1688
rect -1689 712 -1677 1688
rect -1735 700 -1677 712
rect -1477 1688 -1419 1700
rect -1477 712 -1465 1688
rect -1431 712 -1419 1688
rect -1477 700 -1419 712
rect -1319 1688 -1261 1700
rect -1319 712 -1307 1688
rect -1273 712 -1261 1688
rect -1319 700 -1261 712
rect -1061 1688 -1003 1700
rect -1061 712 -1049 1688
rect -1015 712 -1003 1688
rect -1061 700 -1003 712
rect -803 1688 -745 1700
rect -803 712 -791 1688
rect -757 712 -745 1688
rect -803 700 -745 712
rect -545 1688 -487 1700
rect -545 712 -533 1688
rect -499 712 -487 1688
rect -545 700 -487 712
rect -287 1688 -229 1700
rect -287 712 -275 1688
rect -241 712 -229 1688
rect -287 700 -229 712
rect -29 1688 29 1700
rect -29 712 -17 1688
rect 17 712 29 1688
rect -29 700 29 712
rect 229 1688 287 1700
rect 229 712 241 1688
rect 275 712 287 1688
rect 229 700 287 712
rect 487 1688 545 1700
rect 487 712 499 1688
rect 533 712 545 1688
rect 487 700 545 712
rect 745 1688 803 1700
rect 745 712 757 1688
rect 791 712 803 1688
rect 745 700 803 712
rect 1003 1688 1061 1700
rect 1003 712 1015 1688
rect 1049 712 1061 1688
rect 1003 700 1061 712
rect 1261 1688 1319 1700
rect 1261 712 1273 1688
rect 1307 712 1319 1688
rect 1261 700 1319 712
rect 1419 1688 1477 1700
rect 1419 712 1431 1688
rect 1465 712 1477 1688
rect 1419 700 1477 712
rect 1677 1688 1735 1700
rect 1677 712 1689 1688
rect 1723 712 1735 1688
rect 1677 700 1735 712
<< mvndiffc >>
rect -1723 -1688 -1689 -712
rect -1465 -1688 -1431 -712
rect -1307 -1688 -1273 -712
rect -1049 -1688 -1015 -712
rect -791 -1688 -757 -712
rect -533 -1688 -499 -712
rect -275 -1688 -241 -712
rect -17 -1688 17 -712
rect 241 -1688 275 -712
rect 499 -1688 533 -712
rect 757 -1688 791 -712
rect 1015 -1688 1049 -712
rect 1273 -1688 1307 -712
rect 1431 -1688 1465 -712
rect 1689 -1688 1723 -712
rect -2339 -3488 -2305 -2512
rect -2081 -3488 -2047 -2512
rect -1823 -3488 -1789 -2512
rect -1565 -3488 -1531 -2512
rect -1307 -3488 -1273 -2512
rect -1049 -3488 -1015 -2512
rect -791 -3488 -757 -2512
rect -533 -3488 -499 -2512
rect -275 -3488 -241 -2512
rect -17 -3488 17 -2512
rect 241 -3488 275 -2512
rect 499 -3488 533 -2512
rect 757 -3488 791 -2512
rect 1015 -3488 1049 -2512
rect 1273 -3488 1307 -2512
rect 1531 -3488 1565 -2512
rect 1789 -3488 1823 -2512
rect 2047 -3488 2081 -2512
rect 2305 -3488 2339 -2512
<< mvpdiffc >>
rect -2339 2512 -2305 3488
rect -2081 2512 -2047 3488
rect -1823 2512 -1789 3488
rect -1565 2512 -1531 3488
rect -1307 2512 -1273 3488
rect -1049 2512 -1015 3488
rect -791 2512 -757 3488
rect -533 2512 -499 3488
rect -275 2512 -241 3488
rect -17 2512 17 3488
rect 241 2512 275 3488
rect 499 2512 533 3488
rect 757 2512 791 3488
rect 1015 2512 1049 3488
rect 1273 2512 1307 3488
rect 1531 2512 1565 3488
rect 1789 2512 1823 3488
rect 2047 2512 2081 3488
rect 2305 2512 2339 3488
rect -1723 712 -1689 1688
rect -1465 712 -1431 1688
rect -1307 712 -1273 1688
rect -1049 712 -1015 1688
rect -791 712 -757 1688
rect -533 712 -499 1688
rect -275 712 -241 1688
rect -17 712 17 1688
rect 241 712 275 1688
rect 499 712 533 1688
rect 757 712 791 1688
rect 1015 712 1049 1688
rect 1273 712 1307 1688
rect 1431 712 1465 1688
rect 1689 712 1723 1688
<< mvpsubdiff >>
rect -2934 -118 2934 -106
rect -2934 -218 -2760 -118
rect 2760 -218 2934 -118
rect -2934 -230 2934 -218
rect -2934 -280 -2810 -230
rect -2934 -4260 -2922 -280
rect -2822 -4260 -2810 -280
rect 2810 -280 2934 -230
rect -2934 -4310 -2810 -4260
rect 2810 -4260 2822 -280
rect 2922 -4260 2934 -280
rect 2810 -4310 2934 -4260
rect -2934 -4322 2934 -4310
rect -2934 -4422 -2760 -4322
rect 2760 -4422 2934 -4322
rect -2934 -4434 2934 -4422
<< mvnsubdiff >>
rect -2934 4422 2934 4434
rect -2934 4322 -2760 4422
rect 2760 4322 2934 4422
rect -2934 4310 2934 4322
rect -2934 4260 -2810 4310
rect -2934 280 -2922 4260
rect -2822 280 -2810 4260
rect 2810 4260 2934 4310
rect -2934 230 -2810 280
rect 2810 280 2822 4260
rect 2922 280 2934 4260
rect 2810 230 2934 280
rect -2934 218 2934 230
rect -2934 118 -2760 218
rect 2760 118 2934 218
rect -2934 106 2934 118
<< mvpsubdiffcont >>
rect -2760 -218 2760 -118
rect -2922 -4260 -2822 -280
rect 2822 -4260 2922 -280
rect -2760 -4422 2760 -4322
<< mvnsubdiffcont >>
rect -2760 4322 2760 4422
rect -2922 280 -2822 4260
rect 2822 280 2922 4260
rect -2760 118 2760 218
<< poly >>
rect -2259 3581 -2127 3597
rect -2259 3564 -2243 3581
rect -2293 3547 -2243 3564
rect -2143 3564 -2127 3581
rect -2001 3581 -1869 3597
rect -2001 3564 -1985 3581
rect -2143 3547 -2093 3564
rect -2293 3500 -2093 3547
rect -2035 3547 -1985 3564
rect -1885 3564 -1869 3581
rect -1743 3581 -1611 3597
rect -1743 3564 -1727 3581
rect -1885 3547 -1835 3564
rect -2035 3500 -1835 3547
rect -1777 3547 -1727 3564
rect -1627 3564 -1611 3581
rect -1485 3581 -1353 3597
rect -1485 3564 -1469 3581
rect -1627 3547 -1577 3564
rect -1777 3500 -1577 3547
rect -1519 3547 -1469 3564
rect -1369 3564 -1353 3581
rect -1227 3581 -1095 3597
rect -1227 3564 -1211 3581
rect -1369 3547 -1319 3564
rect -1519 3500 -1319 3547
rect -1261 3547 -1211 3564
rect -1111 3564 -1095 3581
rect -969 3581 -837 3597
rect -969 3564 -953 3581
rect -1111 3547 -1061 3564
rect -1261 3500 -1061 3547
rect -1003 3547 -953 3564
rect -853 3564 -837 3581
rect -711 3581 -579 3597
rect -711 3564 -695 3581
rect -853 3547 -803 3564
rect -1003 3500 -803 3547
rect -745 3547 -695 3564
rect -595 3564 -579 3581
rect -453 3581 -321 3597
rect -453 3564 -437 3581
rect -595 3547 -545 3564
rect -745 3500 -545 3547
rect -487 3547 -437 3564
rect -337 3564 -321 3581
rect -195 3581 -63 3597
rect -195 3564 -179 3581
rect -337 3547 -287 3564
rect -487 3500 -287 3547
rect -229 3547 -179 3564
rect -79 3564 -63 3581
rect 63 3581 195 3597
rect 63 3564 79 3581
rect -79 3547 -29 3564
rect -229 3500 -29 3547
rect 29 3547 79 3564
rect 179 3564 195 3581
rect 321 3581 453 3597
rect 321 3564 337 3581
rect 179 3547 229 3564
rect 29 3500 229 3547
rect 287 3547 337 3564
rect 437 3564 453 3581
rect 579 3581 711 3597
rect 579 3564 595 3581
rect 437 3547 487 3564
rect 287 3500 487 3547
rect 545 3547 595 3564
rect 695 3564 711 3581
rect 837 3581 969 3597
rect 837 3564 853 3581
rect 695 3547 745 3564
rect 545 3500 745 3547
rect 803 3547 853 3564
rect 953 3564 969 3581
rect 1095 3581 1227 3597
rect 1095 3564 1111 3581
rect 953 3547 1003 3564
rect 803 3500 1003 3547
rect 1061 3547 1111 3564
rect 1211 3564 1227 3581
rect 1353 3581 1485 3597
rect 1353 3564 1369 3581
rect 1211 3547 1261 3564
rect 1061 3500 1261 3547
rect 1319 3547 1369 3564
rect 1469 3564 1485 3581
rect 1611 3581 1743 3597
rect 1611 3564 1627 3581
rect 1469 3547 1519 3564
rect 1319 3500 1519 3547
rect 1577 3547 1627 3564
rect 1727 3564 1743 3581
rect 1869 3581 2001 3597
rect 1869 3564 1885 3581
rect 1727 3547 1777 3564
rect 1577 3500 1777 3547
rect 1835 3547 1885 3564
rect 1985 3564 2001 3581
rect 2127 3581 2259 3597
rect 2127 3564 2143 3581
rect 1985 3547 2035 3564
rect 1835 3500 2035 3547
rect 2093 3547 2143 3564
rect 2243 3564 2259 3581
rect 2243 3547 2293 3564
rect 2093 3500 2293 3547
rect -2293 2453 -2093 2500
rect -2293 2436 -2243 2453
rect -2259 2419 -2243 2436
rect -2143 2436 -2093 2453
rect -2035 2453 -1835 2500
rect -2035 2436 -1985 2453
rect -2143 2419 -2127 2436
rect -2259 2403 -2127 2419
rect -2001 2419 -1985 2436
rect -1885 2436 -1835 2453
rect -1777 2453 -1577 2500
rect -1777 2436 -1727 2453
rect -1885 2419 -1869 2436
rect -2001 2403 -1869 2419
rect -1743 2419 -1727 2436
rect -1627 2436 -1577 2453
rect -1519 2453 -1319 2500
rect -1519 2436 -1469 2453
rect -1627 2419 -1611 2436
rect -1743 2403 -1611 2419
rect -1485 2419 -1469 2436
rect -1369 2436 -1319 2453
rect -1261 2453 -1061 2500
rect -1261 2436 -1211 2453
rect -1369 2419 -1353 2436
rect -1485 2403 -1353 2419
rect -1227 2419 -1211 2436
rect -1111 2436 -1061 2453
rect -1003 2453 -803 2500
rect -1003 2436 -953 2453
rect -1111 2419 -1095 2436
rect -1227 2403 -1095 2419
rect -969 2419 -953 2436
rect -853 2436 -803 2453
rect -745 2453 -545 2500
rect -745 2436 -695 2453
rect -853 2419 -837 2436
rect -969 2403 -837 2419
rect -711 2419 -695 2436
rect -595 2436 -545 2453
rect -487 2453 -287 2500
rect -487 2436 -437 2453
rect -595 2419 -579 2436
rect -711 2403 -579 2419
rect -453 2419 -437 2436
rect -337 2436 -287 2453
rect -229 2453 -29 2500
rect -229 2436 -179 2453
rect -337 2419 -321 2436
rect -453 2403 -321 2419
rect -195 2419 -179 2436
rect -79 2436 -29 2453
rect 29 2453 229 2500
rect 29 2436 79 2453
rect -79 2419 -63 2436
rect -195 2403 -63 2419
rect 63 2419 79 2436
rect 179 2436 229 2453
rect 287 2453 487 2500
rect 287 2436 337 2453
rect 179 2419 195 2436
rect 63 2403 195 2419
rect 321 2419 337 2436
rect 437 2436 487 2453
rect 545 2453 745 2500
rect 545 2436 595 2453
rect 437 2419 453 2436
rect 321 2403 453 2419
rect 579 2419 595 2436
rect 695 2436 745 2453
rect 803 2453 1003 2500
rect 803 2436 853 2453
rect 695 2419 711 2436
rect 579 2403 711 2419
rect 837 2419 853 2436
rect 953 2436 1003 2453
rect 1061 2453 1261 2500
rect 1061 2436 1111 2453
rect 953 2419 969 2436
rect 837 2403 969 2419
rect 1095 2419 1111 2436
rect 1211 2436 1261 2453
rect 1319 2453 1519 2500
rect 1319 2436 1369 2453
rect 1211 2419 1227 2436
rect 1095 2403 1227 2419
rect 1353 2419 1369 2436
rect 1469 2436 1519 2453
rect 1577 2453 1777 2500
rect 1577 2436 1627 2453
rect 1469 2419 1485 2436
rect 1353 2403 1485 2419
rect 1611 2419 1627 2436
rect 1727 2436 1777 2453
rect 1835 2453 2035 2500
rect 1835 2436 1885 2453
rect 1727 2419 1743 2436
rect 1611 2403 1743 2419
rect 1869 2419 1885 2436
rect 1985 2436 2035 2453
rect 2093 2453 2293 2500
rect 2093 2436 2143 2453
rect 1985 2419 2001 2436
rect 1869 2403 2001 2419
rect 2127 2419 2143 2436
rect 2243 2436 2293 2453
rect 2243 2419 2259 2436
rect 2127 2403 2259 2419
rect -1643 1781 -1511 1797
rect -1643 1764 -1627 1781
rect -1677 1747 -1627 1764
rect -1527 1764 -1511 1781
rect -1419 1781 -1319 1797
rect -1527 1747 -1477 1764
rect -1677 1700 -1477 1747
rect -1419 1747 -1403 1781
rect -1335 1747 -1319 1781
rect -1227 1781 -1095 1797
rect -1227 1764 -1211 1781
rect -1419 1700 -1319 1747
rect -1261 1747 -1211 1764
rect -1111 1764 -1095 1781
rect -969 1781 -837 1797
rect -969 1764 -953 1781
rect -1111 1747 -1061 1764
rect -1261 1700 -1061 1747
rect -1003 1747 -953 1764
rect -853 1764 -837 1781
rect -711 1781 -579 1797
rect -711 1764 -695 1781
rect -853 1747 -803 1764
rect -1003 1700 -803 1747
rect -745 1747 -695 1764
rect -595 1764 -579 1781
rect -453 1781 -321 1797
rect -453 1764 -437 1781
rect -595 1747 -545 1764
rect -745 1700 -545 1747
rect -487 1747 -437 1764
rect -337 1764 -321 1781
rect -195 1781 -63 1797
rect -195 1764 -179 1781
rect -337 1747 -287 1764
rect -487 1700 -287 1747
rect -229 1747 -179 1764
rect -79 1764 -63 1781
rect 63 1781 195 1797
rect 63 1764 79 1781
rect -79 1747 -29 1764
rect -229 1700 -29 1747
rect 29 1747 79 1764
rect 179 1764 195 1781
rect 321 1781 453 1797
rect 321 1764 337 1781
rect 179 1747 229 1764
rect 29 1700 229 1747
rect 287 1747 337 1764
rect 437 1764 453 1781
rect 579 1781 711 1797
rect 579 1764 595 1781
rect 437 1747 487 1764
rect 287 1700 487 1747
rect 545 1747 595 1764
rect 695 1764 711 1781
rect 837 1781 969 1797
rect 837 1764 853 1781
rect 695 1747 745 1764
rect 545 1700 745 1747
rect 803 1747 853 1764
rect 953 1764 969 1781
rect 1095 1781 1227 1797
rect 1095 1764 1111 1781
rect 953 1747 1003 1764
rect 803 1700 1003 1747
rect 1061 1747 1111 1764
rect 1211 1764 1227 1781
rect 1319 1781 1419 1797
rect 1211 1747 1261 1764
rect 1061 1700 1261 1747
rect 1319 1747 1335 1781
rect 1403 1747 1419 1781
rect 1511 1781 1643 1797
rect 1511 1764 1527 1781
rect 1319 1700 1419 1747
rect 1477 1747 1527 1764
rect 1627 1764 1643 1781
rect 1627 1747 1677 1764
rect 1477 1700 1677 1747
rect -1677 653 -1477 700
rect -1677 636 -1627 653
rect -1643 619 -1627 636
rect -1527 636 -1477 653
rect -1419 653 -1319 700
rect -1527 619 -1511 636
rect -1643 603 -1511 619
rect -1419 619 -1403 653
rect -1335 619 -1319 653
rect -1261 653 -1061 700
rect -1261 636 -1211 653
rect -1419 603 -1319 619
rect -1227 619 -1211 636
rect -1111 636 -1061 653
rect -1003 653 -803 700
rect -1003 636 -953 653
rect -1111 619 -1095 636
rect -1227 603 -1095 619
rect -969 619 -953 636
rect -853 636 -803 653
rect -745 653 -545 700
rect -745 636 -695 653
rect -853 619 -837 636
rect -969 603 -837 619
rect -711 619 -695 636
rect -595 636 -545 653
rect -487 653 -287 700
rect -487 636 -437 653
rect -595 619 -579 636
rect -711 603 -579 619
rect -453 619 -437 636
rect -337 636 -287 653
rect -229 653 -29 700
rect -229 636 -179 653
rect -337 619 -321 636
rect -453 603 -321 619
rect -195 619 -179 636
rect -79 636 -29 653
rect 29 653 229 700
rect 29 636 79 653
rect -79 619 -63 636
rect -195 603 -63 619
rect 63 619 79 636
rect 179 636 229 653
rect 287 653 487 700
rect 287 636 337 653
rect 179 619 195 636
rect 63 603 195 619
rect 321 619 337 636
rect 437 636 487 653
rect 545 653 745 700
rect 545 636 595 653
rect 437 619 453 636
rect 321 603 453 619
rect 579 619 595 636
rect 695 636 745 653
rect 803 653 1003 700
rect 803 636 853 653
rect 695 619 711 636
rect 579 603 711 619
rect 837 619 853 636
rect 953 636 1003 653
rect 1061 653 1261 700
rect 1061 636 1111 653
rect 953 619 969 636
rect 837 603 969 619
rect 1095 619 1111 636
rect 1211 636 1261 653
rect 1319 653 1419 700
rect 1211 619 1227 636
rect 1095 603 1227 619
rect 1319 619 1335 653
rect 1403 619 1419 653
rect 1477 653 1677 700
rect 1477 636 1527 653
rect 1319 603 1419 619
rect 1511 619 1527 636
rect 1627 636 1677 653
rect 1627 619 1643 636
rect 1511 603 1643 619
rect -1643 -628 -1511 -612
rect -1643 -645 -1627 -628
rect -1677 -662 -1627 -645
rect -1527 -645 -1511 -628
rect -1419 -628 -1319 -612
rect -1527 -662 -1477 -645
rect -1677 -700 -1477 -662
rect -1419 -662 -1403 -628
rect -1335 -662 -1319 -628
rect -1227 -628 -1095 -612
rect -1227 -645 -1211 -628
rect -1419 -700 -1319 -662
rect -1261 -662 -1211 -645
rect -1111 -645 -1095 -628
rect -969 -628 -837 -612
rect -969 -645 -953 -628
rect -1111 -662 -1061 -645
rect -1261 -700 -1061 -662
rect -1003 -662 -953 -645
rect -853 -645 -837 -628
rect -711 -628 -579 -612
rect -711 -645 -695 -628
rect -853 -662 -803 -645
rect -1003 -700 -803 -662
rect -745 -662 -695 -645
rect -595 -645 -579 -628
rect -453 -628 -321 -612
rect -453 -645 -437 -628
rect -595 -662 -545 -645
rect -745 -700 -545 -662
rect -487 -662 -437 -645
rect -337 -645 -321 -628
rect -195 -628 -63 -612
rect -195 -645 -179 -628
rect -337 -662 -287 -645
rect -487 -700 -287 -662
rect -229 -662 -179 -645
rect -79 -645 -63 -628
rect 63 -628 195 -612
rect 63 -645 79 -628
rect -79 -662 -29 -645
rect -229 -700 -29 -662
rect 29 -662 79 -645
rect 179 -645 195 -628
rect 321 -628 453 -612
rect 321 -645 337 -628
rect 179 -662 229 -645
rect 29 -700 229 -662
rect 287 -662 337 -645
rect 437 -645 453 -628
rect 579 -628 711 -612
rect 579 -645 595 -628
rect 437 -662 487 -645
rect 287 -700 487 -662
rect 545 -662 595 -645
rect 695 -645 711 -628
rect 837 -628 969 -612
rect 837 -645 853 -628
rect 695 -662 745 -645
rect 545 -700 745 -662
rect 803 -662 853 -645
rect 953 -645 969 -628
rect 1095 -628 1227 -612
rect 1095 -645 1111 -628
rect 953 -662 1003 -645
rect 803 -700 1003 -662
rect 1061 -662 1111 -645
rect 1211 -645 1227 -628
rect 1319 -628 1419 -612
rect 1211 -662 1261 -645
rect 1061 -700 1261 -662
rect 1319 -662 1335 -628
rect 1403 -662 1419 -628
rect 1511 -628 1643 -612
rect 1511 -645 1527 -628
rect 1319 -700 1419 -662
rect 1477 -662 1527 -645
rect 1627 -645 1643 -628
rect 1627 -662 1677 -645
rect 1477 -700 1677 -662
rect -1677 -1738 -1477 -1700
rect -1677 -1755 -1627 -1738
rect -1643 -1772 -1627 -1755
rect -1527 -1755 -1477 -1738
rect -1419 -1738 -1319 -1700
rect -1527 -1772 -1511 -1755
rect -1643 -1788 -1511 -1772
rect -1419 -1772 -1403 -1738
rect -1335 -1772 -1319 -1738
rect -1261 -1738 -1061 -1700
rect -1261 -1755 -1211 -1738
rect -1419 -1788 -1319 -1772
rect -1227 -1772 -1211 -1755
rect -1111 -1755 -1061 -1738
rect -1003 -1738 -803 -1700
rect -1003 -1755 -953 -1738
rect -1111 -1772 -1095 -1755
rect -1227 -1788 -1095 -1772
rect -969 -1772 -953 -1755
rect -853 -1755 -803 -1738
rect -745 -1738 -545 -1700
rect -745 -1755 -695 -1738
rect -853 -1772 -837 -1755
rect -969 -1788 -837 -1772
rect -711 -1772 -695 -1755
rect -595 -1755 -545 -1738
rect -487 -1738 -287 -1700
rect -487 -1755 -437 -1738
rect -595 -1772 -579 -1755
rect -711 -1788 -579 -1772
rect -453 -1772 -437 -1755
rect -337 -1755 -287 -1738
rect -229 -1738 -29 -1700
rect -229 -1755 -179 -1738
rect -337 -1772 -321 -1755
rect -453 -1788 -321 -1772
rect -195 -1772 -179 -1755
rect -79 -1755 -29 -1738
rect 29 -1738 229 -1700
rect 29 -1755 79 -1738
rect -79 -1772 -63 -1755
rect -195 -1788 -63 -1772
rect 63 -1772 79 -1755
rect 179 -1755 229 -1738
rect 287 -1738 487 -1700
rect 287 -1755 337 -1738
rect 179 -1772 195 -1755
rect 63 -1788 195 -1772
rect 321 -1772 337 -1755
rect 437 -1755 487 -1738
rect 545 -1738 745 -1700
rect 545 -1755 595 -1738
rect 437 -1772 453 -1755
rect 321 -1788 453 -1772
rect 579 -1772 595 -1755
rect 695 -1755 745 -1738
rect 803 -1738 1003 -1700
rect 803 -1755 853 -1738
rect 695 -1772 711 -1755
rect 579 -1788 711 -1772
rect 837 -1772 853 -1755
rect 953 -1755 1003 -1738
rect 1061 -1738 1261 -1700
rect 1061 -1755 1111 -1738
rect 953 -1772 969 -1755
rect 837 -1788 969 -1772
rect 1095 -1772 1111 -1755
rect 1211 -1755 1261 -1738
rect 1319 -1738 1419 -1700
rect 1211 -1772 1227 -1755
rect 1095 -1788 1227 -1772
rect 1319 -1772 1335 -1738
rect 1403 -1772 1419 -1738
rect 1477 -1738 1677 -1700
rect 1477 -1755 1527 -1738
rect 1319 -1788 1419 -1772
rect 1511 -1772 1527 -1755
rect 1627 -1755 1677 -1738
rect 1627 -1772 1643 -1755
rect 1511 -1788 1643 -1772
rect -2259 -2428 -2127 -2412
rect -2259 -2445 -2243 -2428
rect -2293 -2462 -2243 -2445
rect -2143 -2445 -2127 -2428
rect -2001 -2428 -1869 -2412
rect -2001 -2445 -1985 -2428
rect -2143 -2462 -2093 -2445
rect -2293 -2500 -2093 -2462
rect -2035 -2462 -1985 -2445
rect -1885 -2445 -1869 -2428
rect -1743 -2428 -1611 -2412
rect -1743 -2445 -1727 -2428
rect -1885 -2462 -1835 -2445
rect -2035 -2500 -1835 -2462
rect -1777 -2462 -1727 -2445
rect -1627 -2445 -1611 -2428
rect -1485 -2428 -1353 -2412
rect -1485 -2445 -1469 -2428
rect -1627 -2462 -1577 -2445
rect -1777 -2500 -1577 -2462
rect -1519 -2462 -1469 -2445
rect -1369 -2445 -1353 -2428
rect -1227 -2428 -1095 -2412
rect -1227 -2445 -1211 -2428
rect -1369 -2462 -1319 -2445
rect -1519 -2500 -1319 -2462
rect -1261 -2462 -1211 -2445
rect -1111 -2445 -1095 -2428
rect -969 -2428 -837 -2412
rect -969 -2445 -953 -2428
rect -1111 -2462 -1061 -2445
rect -1261 -2500 -1061 -2462
rect -1003 -2462 -953 -2445
rect -853 -2445 -837 -2428
rect -711 -2428 -579 -2412
rect -711 -2445 -695 -2428
rect -853 -2462 -803 -2445
rect -1003 -2500 -803 -2462
rect -745 -2462 -695 -2445
rect -595 -2445 -579 -2428
rect -453 -2428 -321 -2412
rect -453 -2445 -437 -2428
rect -595 -2462 -545 -2445
rect -745 -2500 -545 -2462
rect -487 -2462 -437 -2445
rect -337 -2445 -321 -2428
rect -195 -2428 -63 -2412
rect -195 -2445 -179 -2428
rect -337 -2462 -287 -2445
rect -487 -2500 -287 -2462
rect -229 -2462 -179 -2445
rect -79 -2445 -63 -2428
rect 63 -2428 195 -2412
rect 63 -2445 79 -2428
rect -79 -2462 -29 -2445
rect -229 -2500 -29 -2462
rect 29 -2462 79 -2445
rect 179 -2445 195 -2428
rect 321 -2428 453 -2412
rect 321 -2445 337 -2428
rect 179 -2462 229 -2445
rect 29 -2500 229 -2462
rect 287 -2462 337 -2445
rect 437 -2445 453 -2428
rect 579 -2428 711 -2412
rect 579 -2445 595 -2428
rect 437 -2462 487 -2445
rect 287 -2500 487 -2462
rect 545 -2462 595 -2445
rect 695 -2445 711 -2428
rect 837 -2428 969 -2412
rect 837 -2445 853 -2428
rect 695 -2462 745 -2445
rect 545 -2500 745 -2462
rect 803 -2462 853 -2445
rect 953 -2445 969 -2428
rect 1095 -2428 1227 -2412
rect 1095 -2445 1111 -2428
rect 953 -2462 1003 -2445
rect 803 -2500 1003 -2462
rect 1061 -2462 1111 -2445
rect 1211 -2445 1227 -2428
rect 1353 -2428 1485 -2412
rect 1353 -2445 1369 -2428
rect 1211 -2462 1261 -2445
rect 1061 -2500 1261 -2462
rect 1319 -2462 1369 -2445
rect 1469 -2445 1485 -2428
rect 1611 -2428 1743 -2412
rect 1611 -2445 1627 -2428
rect 1469 -2462 1519 -2445
rect 1319 -2500 1519 -2462
rect 1577 -2462 1627 -2445
rect 1727 -2445 1743 -2428
rect 1869 -2428 2001 -2412
rect 1869 -2445 1885 -2428
rect 1727 -2462 1777 -2445
rect 1577 -2500 1777 -2462
rect 1835 -2462 1885 -2445
rect 1985 -2445 2001 -2428
rect 2127 -2428 2259 -2412
rect 2127 -2445 2143 -2428
rect 1985 -2462 2035 -2445
rect 1835 -2500 2035 -2462
rect 2093 -2462 2143 -2445
rect 2243 -2445 2259 -2428
rect 2243 -2462 2293 -2445
rect 2093 -2500 2293 -2462
rect -2293 -3538 -2093 -3500
rect -2293 -3555 -2243 -3538
rect -2259 -3572 -2243 -3555
rect -2143 -3555 -2093 -3538
rect -2035 -3538 -1835 -3500
rect -2035 -3555 -1985 -3538
rect -2143 -3572 -2127 -3555
rect -2259 -3588 -2127 -3572
rect -2001 -3572 -1985 -3555
rect -1885 -3555 -1835 -3538
rect -1777 -3538 -1577 -3500
rect -1777 -3555 -1727 -3538
rect -1885 -3572 -1869 -3555
rect -2001 -3588 -1869 -3572
rect -1743 -3572 -1727 -3555
rect -1627 -3555 -1577 -3538
rect -1519 -3538 -1319 -3500
rect -1519 -3555 -1469 -3538
rect -1627 -3572 -1611 -3555
rect -1743 -3588 -1611 -3572
rect -1485 -3572 -1469 -3555
rect -1369 -3555 -1319 -3538
rect -1261 -3538 -1061 -3500
rect -1261 -3555 -1211 -3538
rect -1369 -3572 -1353 -3555
rect -1485 -3588 -1353 -3572
rect -1227 -3572 -1211 -3555
rect -1111 -3555 -1061 -3538
rect -1003 -3538 -803 -3500
rect -1003 -3555 -953 -3538
rect -1111 -3572 -1095 -3555
rect -1227 -3588 -1095 -3572
rect -969 -3572 -953 -3555
rect -853 -3555 -803 -3538
rect -745 -3538 -545 -3500
rect -745 -3555 -695 -3538
rect -853 -3572 -837 -3555
rect -969 -3588 -837 -3572
rect -711 -3572 -695 -3555
rect -595 -3555 -545 -3538
rect -487 -3538 -287 -3500
rect -487 -3555 -437 -3538
rect -595 -3572 -579 -3555
rect -711 -3588 -579 -3572
rect -453 -3572 -437 -3555
rect -337 -3555 -287 -3538
rect -229 -3538 -29 -3500
rect -229 -3555 -179 -3538
rect -337 -3572 -321 -3555
rect -453 -3588 -321 -3572
rect -195 -3572 -179 -3555
rect -79 -3555 -29 -3538
rect 29 -3538 229 -3500
rect 29 -3555 79 -3538
rect -79 -3572 -63 -3555
rect -195 -3588 -63 -3572
rect 63 -3572 79 -3555
rect 179 -3555 229 -3538
rect 287 -3538 487 -3500
rect 287 -3555 337 -3538
rect 179 -3572 195 -3555
rect 63 -3588 195 -3572
rect 321 -3572 337 -3555
rect 437 -3555 487 -3538
rect 545 -3538 745 -3500
rect 545 -3555 595 -3538
rect 437 -3572 453 -3555
rect 321 -3588 453 -3572
rect 579 -3572 595 -3555
rect 695 -3555 745 -3538
rect 803 -3538 1003 -3500
rect 803 -3555 853 -3538
rect 695 -3572 711 -3555
rect 579 -3588 711 -3572
rect 837 -3572 853 -3555
rect 953 -3555 1003 -3538
rect 1061 -3538 1261 -3500
rect 1061 -3555 1111 -3538
rect 953 -3572 969 -3555
rect 837 -3588 969 -3572
rect 1095 -3572 1111 -3555
rect 1211 -3555 1261 -3538
rect 1319 -3538 1519 -3500
rect 1319 -3555 1369 -3538
rect 1211 -3572 1227 -3555
rect 1095 -3588 1227 -3572
rect 1353 -3572 1369 -3555
rect 1469 -3555 1519 -3538
rect 1577 -3538 1777 -3500
rect 1577 -3555 1627 -3538
rect 1469 -3572 1485 -3555
rect 1353 -3588 1485 -3572
rect 1611 -3572 1627 -3555
rect 1727 -3555 1777 -3538
rect 1835 -3538 2035 -3500
rect 1835 -3555 1885 -3538
rect 1727 -3572 1743 -3555
rect 1611 -3588 1743 -3572
rect 1869 -3572 1885 -3555
rect 1985 -3555 2035 -3538
rect 2093 -3538 2293 -3500
rect 2093 -3555 2143 -3538
rect 1985 -3572 2001 -3555
rect 1869 -3588 2001 -3572
rect 2127 -3572 2143 -3555
rect 2243 -3555 2293 -3538
rect 2243 -3572 2259 -3555
rect 2127 -3588 2259 -3572
<< polycont >>
rect -2243 3547 -2143 3581
rect -1985 3547 -1885 3581
rect -1727 3547 -1627 3581
rect -1469 3547 -1369 3581
rect -1211 3547 -1111 3581
rect -953 3547 -853 3581
rect -695 3547 -595 3581
rect -437 3547 -337 3581
rect -179 3547 -79 3581
rect 79 3547 179 3581
rect 337 3547 437 3581
rect 595 3547 695 3581
rect 853 3547 953 3581
rect 1111 3547 1211 3581
rect 1369 3547 1469 3581
rect 1627 3547 1727 3581
rect 1885 3547 1985 3581
rect 2143 3547 2243 3581
rect -2243 2419 -2143 2453
rect -1985 2419 -1885 2453
rect -1727 2419 -1627 2453
rect -1469 2419 -1369 2453
rect -1211 2419 -1111 2453
rect -953 2419 -853 2453
rect -695 2419 -595 2453
rect -437 2419 -337 2453
rect -179 2419 -79 2453
rect 79 2419 179 2453
rect 337 2419 437 2453
rect 595 2419 695 2453
rect 853 2419 953 2453
rect 1111 2419 1211 2453
rect 1369 2419 1469 2453
rect 1627 2419 1727 2453
rect 1885 2419 1985 2453
rect 2143 2419 2243 2453
rect -1627 1747 -1527 1781
rect -1403 1747 -1335 1781
rect -1211 1747 -1111 1781
rect -953 1747 -853 1781
rect -695 1747 -595 1781
rect -437 1747 -337 1781
rect -179 1747 -79 1781
rect 79 1747 179 1781
rect 337 1747 437 1781
rect 595 1747 695 1781
rect 853 1747 953 1781
rect 1111 1747 1211 1781
rect 1335 1747 1403 1781
rect 1527 1747 1627 1781
rect -1627 619 -1527 653
rect -1403 619 -1335 653
rect -1211 619 -1111 653
rect -953 619 -853 653
rect -695 619 -595 653
rect -437 619 -337 653
rect -179 619 -79 653
rect 79 619 179 653
rect 337 619 437 653
rect 595 619 695 653
rect 853 619 953 653
rect 1111 619 1211 653
rect 1335 619 1403 653
rect 1527 619 1627 653
rect -1627 -662 -1527 -628
rect -1403 -662 -1335 -628
rect -1211 -662 -1111 -628
rect -953 -662 -853 -628
rect -695 -662 -595 -628
rect -437 -662 -337 -628
rect -179 -662 -79 -628
rect 79 -662 179 -628
rect 337 -662 437 -628
rect 595 -662 695 -628
rect 853 -662 953 -628
rect 1111 -662 1211 -628
rect 1335 -662 1403 -628
rect 1527 -662 1627 -628
rect -1627 -1772 -1527 -1738
rect -1403 -1772 -1335 -1738
rect -1211 -1772 -1111 -1738
rect -953 -1772 -853 -1738
rect -695 -1772 -595 -1738
rect -437 -1772 -337 -1738
rect -179 -1772 -79 -1738
rect 79 -1772 179 -1738
rect 337 -1772 437 -1738
rect 595 -1772 695 -1738
rect 853 -1772 953 -1738
rect 1111 -1772 1211 -1738
rect 1335 -1772 1403 -1738
rect 1527 -1772 1627 -1738
rect -2243 -2462 -2143 -2428
rect -1985 -2462 -1885 -2428
rect -1727 -2462 -1627 -2428
rect -1469 -2462 -1369 -2428
rect -1211 -2462 -1111 -2428
rect -953 -2462 -853 -2428
rect -695 -2462 -595 -2428
rect -437 -2462 -337 -2428
rect -179 -2462 -79 -2428
rect 79 -2462 179 -2428
rect 337 -2462 437 -2428
rect 595 -2462 695 -2428
rect 853 -2462 953 -2428
rect 1111 -2462 1211 -2428
rect 1369 -2462 1469 -2428
rect 1627 -2462 1727 -2428
rect 1885 -2462 1985 -2428
rect 2143 -2462 2243 -2428
rect -2243 -3572 -2143 -3538
rect -1985 -3572 -1885 -3538
rect -1727 -3572 -1627 -3538
rect -1469 -3572 -1369 -3538
rect -1211 -3572 -1111 -3538
rect -953 -3572 -853 -3538
rect -695 -3572 -595 -3538
rect -437 -3572 -337 -3538
rect -179 -3572 -79 -3538
rect 79 -3572 179 -3538
rect 337 -3572 437 -3538
rect 595 -3572 695 -3538
rect 853 -3572 953 -3538
rect 1111 -3572 1211 -3538
rect 1369 -3572 1469 -3538
rect 1627 -3572 1727 -3538
rect 1885 -3572 1985 -3538
rect 2143 -3572 2243 -3538
<< locali >>
rect -2922 4260 -2822 4422
rect 2822 4260 2922 4422
rect -2001 3797 2001 4197
rect -2001 3581 -1869 3797
rect -2259 3547 -2243 3581
rect -2143 3547 -2127 3581
rect -2001 3547 -1985 3581
rect -1885 3547 -1869 3581
rect -1743 3581 -1611 3797
rect -1743 3547 -1727 3581
rect -1627 3547 -1611 3581
rect -1485 3581 -1353 3797
rect -969 3581 -837 3797
rect -1485 3547 -1469 3581
rect -1369 3547 -1353 3581
rect -1227 3547 -1211 3581
rect -1111 3547 -1095 3581
rect -969 3547 -953 3581
rect -853 3547 -837 3581
rect -711 3621 711 3763
rect -711 3581 -579 3621
rect -711 3547 -695 3581
rect -595 3547 -579 3581
rect -453 3581 -321 3621
rect -453 3547 -437 3581
rect -337 3547 -321 3581
rect -195 3581 -63 3621
rect -195 3547 -179 3581
rect -79 3547 -63 3581
rect 62 3581 195 3621
rect 62 3547 79 3581
rect 179 3547 195 3581
rect 321 3581 453 3621
rect 321 3547 337 3581
rect 437 3547 453 3581
rect 579 3581 711 3621
rect 579 3547 595 3581
rect 695 3547 711 3581
rect 837 3581 969 3797
rect 1353 3581 1485 3797
rect 837 3547 853 3581
rect 953 3547 969 3581
rect 1095 3547 1111 3581
rect 1211 3547 1227 3581
rect 1353 3547 1369 3581
rect 1469 3547 1485 3581
rect 1611 3581 1743 3797
rect 1611 3547 1627 3581
rect 1727 3547 1743 3581
rect 1869 3581 2001 3797
rect 1869 3547 1885 3581
rect 1985 3547 2001 3581
rect 2127 3547 2143 3581
rect 2243 3547 2259 3581
rect -2339 3488 -2305 3504
rect -2339 2496 -2305 2512
rect -2081 3488 -2047 3504
rect -2081 2496 -2047 2512
rect -1823 3488 -1789 3504
rect -1823 2496 -1789 2512
rect -1565 3488 -1531 3504
rect -1565 2496 -1531 2512
rect -1307 3488 -1273 3504
rect -1307 2496 -1273 2512
rect -1049 3488 -1015 3504
rect -1049 2496 -1015 2512
rect -791 3488 -757 3504
rect -791 2496 -757 2512
rect -533 3488 -499 3504
rect -533 2496 -499 2512
rect -275 3488 -241 3504
rect -275 2496 -241 2512
rect -17 3488 17 3504
rect -17 2496 17 2512
rect 241 3488 275 3504
rect 241 2496 275 2512
rect 499 3488 533 3504
rect 499 2496 533 2512
rect 757 3488 791 3504
rect 757 2496 791 2512
rect 1015 3488 1049 3504
rect 1015 2496 1049 2512
rect 1273 3488 1307 3504
rect 1273 2496 1307 2512
rect 1531 3488 1565 3504
rect 1531 2496 1565 2512
rect 1789 3488 1823 3504
rect 1789 2496 1823 2512
rect 2047 3488 2081 3504
rect 2047 2496 2081 2512
rect 2305 3488 2339 3504
rect 2305 2496 2339 2512
rect -2259 2419 -2243 2453
rect -2143 2419 -2127 2453
rect -2001 2419 -1985 2453
rect -1885 2419 -1869 2453
rect -1743 2419 -1727 2453
rect -1627 2419 -1611 2453
rect -1485 2419 -1469 2453
rect -1369 2419 -1353 2453
rect -1227 2419 -1211 2453
rect -1111 2419 -1095 2453
rect -969 2419 -953 2453
rect -853 2419 -837 2453
rect -711 2419 -695 2453
rect -595 2419 -579 2453
rect -453 2419 -437 2453
rect -337 2419 -321 2453
rect -195 2419 -179 2453
rect -79 2419 -63 2453
rect 63 2419 79 2453
rect 179 2419 195 2453
rect 321 2419 337 2453
rect 437 2419 453 2453
rect 579 2419 595 2453
rect 695 2419 711 2453
rect 837 2419 853 2453
rect 953 2419 969 2453
rect 1095 2419 1111 2453
rect 1211 2419 1227 2453
rect 1353 2419 1369 2453
rect 1469 2419 1485 2453
rect 1611 2419 1627 2453
rect 1727 2419 1743 2453
rect 1869 2419 1885 2453
rect 1985 2419 2001 2453
rect 2127 2419 2143 2453
rect 2243 2419 2259 2453
rect -1419 2282 1419 2333
rect -1419 2202 -659 2282
rect -579 2202 579 2282
rect 659 2202 1419 2282
rect -1419 2049 1419 2202
rect -1419 1781 -1319 2049
rect -969 2008 969 2015
rect -969 1958 -963 2008
rect -913 1958 913 2008
rect 963 1958 969 2008
rect -969 1821 969 1958
rect -969 1781 -837 1821
rect -195 1781 -63 1821
rect -1643 1747 -1627 1781
rect -1527 1747 -1511 1781
rect -1419 1747 -1403 1781
rect -1335 1747 -1319 1781
rect -1227 1747 -1211 1781
rect -1111 1747 -1095 1781
rect -969 1747 -953 1781
rect -853 1747 -837 1781
rect -711 1747 -695 1781
rect -595 1747 -579 1781
rect -453 1747 -437 1781
rect -337 1747 -321 1781
rect -195 1747 -179 1781
rect -79 1747 -63 1781
rect 63 1781 195 1821
rect 837 1781 969 1821
rect 1319 1781 1419 2049
rect 63 1747 79 1781
rect 179 1747 195 1781
rect 321 1747 337 1781
rect 437 1747 453 1781
rect 579 1747 595 1781
rect 695 1747 711 1781
rect 837 1747 853 1781
rect 953 1747 969 1781
rect 1095 1747 1111 1781
rect 1211 1747 1227 1781
rect 1319 1747 1335 1781
rect 1403 1747 1419 1781
rect 1511 1747 1527 1781
rect 1627 1747 1643 1781
rect -1723 1688 -1689 1704
rect -1723 696 -1689 712
rect -1465 1688 -1431 1704
rect -1465 696 -1431 712
rect -1307 1688 -1273 1704
rect -1307 696 -1273 712
rect -1049 1688 -1015 1704
rect -1049 696 -1015 712
rect -791 1688 -757 1704
rect -791 696 -757 712
rect -533 1688 -499 1704
rect -533 696 -499 712
rect -275 1688 -241 1704
rect -275 696 -241 712
rect -17 1688 17 1704
rect -17 696 17 712
rect 241 1688 275 1704
rect 241 696 275 712
rect 499 1688 533 1704
rect 499 696 533 712
rect 757 1688 791 1704
rect 757 696 791 712
rect 1015 1688 1049 1704
rect 1015 696 1049 712
rect 1273 1688 1307 1704
rect 1273 696 1307 712
rect 1431 1688 1465 1704
rect 1431 696 1465 712
rect 1689 1688 1723 1704
rect 1689 696 1723 712
rect -1643 619 -1627 653
rect -1527 619 -1511 653
rect -1419 619 -1403 653
rect -1335 619 -1319 653
rect -1227 619 -1211 653
rect -1111 619 -1095 653
rect -969 619 -953 653
rect -853 619 -837 653
rect -711 619 -695 653
rect -595 619 -579 653
rect -711 579 -579 619
rect -453 619 -437 653
rect -337 619 -321 653
rect -195 619 -179 653
rect -79 619 -63 653
rect 63 619 79 653
rect 179 619 195 653
rect 321 619 337 653
rect 437 619 453 653
rect -453 579 -321 619
rect 321 579 453 619
rect 579 619 595 653
rect 695 619 711 653
rect 837 619 853 653
rect 953 619 969 653
rect 1095 619 1111 653
rect 1211 619 1227 653
rect 1319 619 1335 653
rect 1403 619 1419 653
rect 1511 619 1527 653
rect 1627 619 1643 653
rect 579 579 711 619
rect -1262 567 1264 579
rect -1212 517 1202 567
rect 1252 517 1264 567
rect -1262 437 1264 517
rect -447 436 -315 437
rect -2922 118 -2822 280
rect 2822 118 2922 280
rect -2922 -280 -2822 -118
rect 2822 -280 2922 -118
rect -969 -458 969 -394
rect -969 -538 -41 -458
rect 39 -538 969 -458
rect -969 -588 969 -538
rect -969 -628 -837 -588
rect -195 -628 -63 -588
rect -1643 -662 -1627 -628
rect -1527 -662 -1511 -628
rect -1419 -662 -1403 -628
rect -1335 -662 -1319 -628
rect -1227 -662 -1211 -628
rect -1111 -662 -1095 -628
rect -969 -662 -953 -628
rect -853 -662 -837 -628
rect -711 -662 -695 -628
rect -595 -662 -579 -628
rect -453 -662 -437 -628
rect -337 -662 -321 -628
rect -195 -662 -179 -628
rect -79 -662 -63 -628
rect 63 -628 195 -588
rect 837 -628 969 -588
rect 63 -662 79 -628
rect 179 -662 195 -628
rect 321 -662 337 -628
rect 437 -662 453 -628
rect 579 -662 595 -628
rect 695 -662 711 -628
rect 837 -662 853 -628
rect 953 -662 969 -628
rect 1095 -662 1111 -628
rect 1211 -662 1227 -628
rect 1319 -662 1335 -628
rect 1403 -662 1419 -628
rect 1511 -662 1527 -628
rect 1627 -662 1643 -628
rect -1723 -712 -1689 -696
rect -1723 -1704 -1689 -1688
rect -1465 -712 -1431 -696
rect -1465 -1704 -1431 -1688
rect -1307 -712 -1273 -696
rect -1307 -1704 -1273 -1688
rect -1049 -712 -1015 -696
rect -1049 -1704 -1015 -1688
rect -791 -712 -757 -696
rect -791 -1704 -757 -1688
rect -533 -712 -499 -696
rect -533 -1704 -499 -1688
rect -275 -712 -241 -696
rect -275 -1704 -241 -1688
rect -17 -712 17 -696
rect -17 -1704 17 -1688
rect 241 -712 275 -696
rect 241 -1704 275 -1688
rect 499 -712 533 -696
rect 499 -1704 533 -1688
rect 757 -712 791 -696
rect 757 -1704 791 -1688
rect 1015 -712 1049 -696
rect 1015 -1704 1049 -1688
rect 1273 -712 1307 -696
rect 1273 -1704 1307 -1688
rect 1431 -712 1465 -696
rect 1431 -1704 1465 -1688
rect 1689 -712 1723 -696
rect 1689 -1704 1723 -1688
rect -1643 -1772 -1627 -1738
rect -1527 -1772 -1511 -1738
rect -1419 -1772 -1403 -1738
rect -1335 -1772 -1319 -1738
rect -1227 -1772 -1211 -1738
rect -1111 -1772 -1095 -1738
rect -969 -1772 -953 -1738
rect -853 -1772 -837 -1738
rect -711 -1772 -695 -1738
rect -595 -1772 -579 -1738
rect -1419 -1988 -1319 -1772
rect -711 -1812 -579 -1772
rect -453 -1772 -437 -1738
rect -337 -1772 -321 -1738
rect -195 -1772 -179 -1738
rect -79 -1772 -63 -1738
rect 63 -1772 79 -1738
rect 179 -1772 195 -1738
rect 321 -1772 337 -1738
rect 437 -1772 453 -1738
rect -453 -1812 -321 -1772
rect 321 -1812 453 -1772
rect 579 -1772 595 -1738
rect 695 -1772 711 -1738
rect 837 -1772 853 -1738
rect 953 -1772 969 -1738
rect 1095 -1772 1111 -1738
rect 1211 -1772 1227 -1738
rect 1319 -1772 1335 -1738
rect 1403 -1772 1419 -1738
rect 1511 -1772 1527 -1738
rect 1627 -1772 1643 -1738
rect 579 -1812 711 -1772
rect -711 -1822 711 -1812
rect -711 -1902 -685 -1822
rect -605 -1902 -427 -1822
rect -347 -1902 347 -1822
rect 427 -1902 605 -1822
rect 685 -1902 711 -1822
rect -711 -1954 711 -1902
rect 1319 -1988 1419 -1772
rect -1419 -2046 1419 -1988
rect -1419 -2126 -556 -2046
rect -476 -2126 476 -2046
rect 556 -2126 1419 -2046
rect -1419 -2272 1419 -2126
rect -2259 -2462 -2243 -2428
rect -2143 -2462 -2127 -2428
rect -2001 -2462 -1985 -2428
rect -1885 -2462 -1869 -2428
rect -1743 -2462 -1727 -2428
rect -1627 -2462 -1611 -2428
rect -1485 -2462 -1469 -2428
rect -1369 -2462 -1353 -2428
rect -1227 -2462 -1211 -2428
rect -1111 -2462 -1095 -2428
rect -969 -2462 -953 -2428
rect -853 -2462 -837 -2428
rect -711 -2462 -695 -2428
rect -595 -2462 -579 -2428
rect -453 -2462 -437 -2428
rect -337 -2462 -321 -2428
rect -195 -2462 -179 -2428
rect -79 -2462 -63 -2428
rect 63 -2462 79 -2428
rect 179 -2462 195 -2428
rect 321 -2462 337 -2428
rect 437 -2462 453 -2428
rect 579 -2462 595 -2428
rect 695 -2462 711 -2428
rect 837 -2462 853 -2428
rect 953 -2462 969 -2428
rect 1095 -2462 1111 -2428
rect 1211 -2462 1227 -2428
rect 1353 -2462 1369 -2428
rect 1469 -2462 1485 -2428
rect 1611 -2462 1627 -2428
rect 1727 -2462 1743 -2428
rect 1869 -2462 1885 -2428
rect 1985 -2462 2001 -2428
rect 2127 -2462 2143 -2428
rect 2243 -2462 2259 -2428
rect -2339 -2512 -2305 -2496
rect -2339 -3504 -2305 -3488
rect -2081 -2512 -2047 -2496
rect -2081 -3504 -2047 -3488
rect -1823 -2512 -1789 -2496
rect -1823 -3504 -1789 -3488
rect -1565 -2512 -1531 -2496
rect -1565 -3504 -1531 -3488
rect -1307 -2512 -1273 -2496
rect -1307 -3504 -1273 -3488
rect -1049 -2512 -1015 -2496
rect -1049 -3504 -1015 -3488
rect -791 -2512 -757 -2496
rect -791 -3504 -757 -3488
rect -533 -2512 -499 -2496
rect -533 -3504 -499 -3488
rect -275 -2512 -241 -2496
rect -275 -3504 -241 -3488
rect -17 -2512 17 -2496
rect -17 -3504 17 -3488
rect 241 -2512 275 -2496
rect 241 -3504 275 -3488
rect 499 -2512 533 -2496
rect 499 -3504 533 -3488
rect 757 -2512 791 -2496
rect 757 -3504 791 -3488
rect 1015 -2512 1049 -2496
rect 1015 -3504 1049 -3488
rect 1273 -2512 1307 -2496
rect 1273 -3504 1307 -3488
rect 1531 -2512 1565 -2496
rect 1531 -3504 1565 -3488
rect 1789 -2512 1823 -2496
rect 1789 -3504 1823 -3488
rect 2047 -2512 2081 -2496
rect 2047 -3504 2081 -3488
rect 2305 -2512 2339 -2496
rect 2305 -3504 2339 -3488
rect -2259 -3572 -2243 -3538
rect -2143 -3572 -2127 -3538
rect -2001 -3572 -1985 -3538
rect -1885 -3572 -1869 -3538
rect -1743 -3572 -1727 -3538
rect -1627 -3572 -1611 -3538
rect -1485 -3572 -1469 -3538
rect -1369 -3572 -1353 -3538
rect -1227 -3572 -1211 -3538
rect -1111 -3572 -1095 -3538
rect -969 -3572 -953 -3538
rect -853 -3572 -837 -3538
rect -711 -3572 -695 -3538
rect -595 -3572 -579 -3538
rect -453 -3572 -437 -3538
rect -337 -3572 -321 -3538
rect -195 -3572 -179 -3538
rect -79 -3572 -63 -3538
rect 63 -3572 79 -3538
rect 179 -3572 195 -3538
rect 321 -3572 337 -3538
rect 437 -3572 453 -3538
rect 579 -3572 595 -3538
rect 695 -3572 711 -3538
rect 837 -3572 853 -3538
rect 953 -3572 969 -3538
rect 1095 -3572 1111 -3538
rect 1211 -3572 1227 -3538
rect 1353 -3572 1369 -3538
rect 1469 -3572 1485 -3538
rect 1611 -3572 1627 -3538
rect 1727 -3572 1743 -3538
rect 1869 -3572 1885 -3538
rect 1985 -3572 2001 -3538
rect 2127 -3572 2143 -3538
rect 2243 -3572 2259 -3538
rect -2922 -4422 -2822 -4260
rect 2822 -4422 2922 -4260
<< viali >>
rect -2822 4322 -2760 4422
rect -2760 4322 2760 4422
rect 2760 4322 2822 4422
rect -2922 423 -2822 4117
rect -2227 3547 -2159 3581
rect -1969 3547 -1901 3581
rect -1711 3547 -1643 3581
rect -1453 3547 -1385 3581
rect -1195 3547 -1127 3581
rect -937 3547 -869 3581
rect -679 3547 -611 3581
rect -421 3547 -353 3581
rect -163 3547 -95 3581
rect 95 3547 163 3581
rect 353 3547 421 3581
rect 611 3547 679 3581
rect 869 3547 937 3581
rect 1127 3547 1195 3581
rect 1385 3547 1453 3581
rect 1643 3547 1711 3581
rect 1901 3547 1969 3581
rect 2159 3547 2227 3581
rect -2339 2512 -2305 3488
rect -2081 2512 -2047 3488
rect -1823 2512 -1789 3488
rect -1565 2512 -1531 3488
rect -1307 2512 -1273 3488
rect -1049 2512 -1015 3488
rect -791 2512 -757 3488
rect -533 2512 -499 3488
rect -275 2512 -241 3488
rect -17 2512 17 3488
rect 241 2512 275 3488
rect 499 2512 533 3488
rect 757 2512 791 3488
rect 1015 2512 1049 3488
rect 1273 2512 1307 3488
rect 1531 2512 1565 3488
rect 1789 2512 1823 3488
rect 2047 2512 2081 3488
rect 2305 2512 2339 3488
rect -2227 2419 -2159 2453
rect -1969 2419 -1901 2453
rect -1711 2419 -1643 2453
rect -1453 2419 -1385 2453
rect -1195 2419 -1127 2453
rect -937 2419 -869 2453
rect -679 2419 -611 2453
rect -421 2419 -353 2453
rect -163 2419 -95 2453
rect 95 2419 163 2453
rect 353 2419 421 2453
rect 611 2419 679 2453
rect 869 2419 937 2453
rect 1127 2419 1195 2453
rect 1385 2419 1453 2453
rect 1643 2419 1711 2453
rect 1901 2419 1969 2453
rect 2159 2419 2227 2453
rect -659 2202 -579 2282
rect 579 2202 659 2282
rect -963 1958 -913 2008
rect 913 1958 963 2008
rect -1611 1747 -1543 1781
rect -1396 1747 -1342 1781
rect -1195 1747 -1127 1781
rect -937 1747 -869 1781
rect -679 1747 -611 1781
rect -421 1747 -353 1781
rect -163 1747 -95 1781
rect 95 1747 163 1781
rect 353 1747 421 1781
rect 611 1747 679 1781
rect 869 1747 937 1781
rect 1127 1747 1195 1781
rect 1342 1747 1396 1781
rect 1543 1747 1611 1781
rect -1723 712 -1689 1688
rect -1465 712 -1431 1688
rect -1307 712 -1273 1688
rect -1049 712 -1015 1688
rect -791 712 -757 1688
rect -533 712 -499 1688
rect -275 712 -241 1688
rect -17 712 17 1688
rect 241 712 275 1688
rect 499 712 533 1688
rect 757 712 791 1688
rect 1015 712 1049 1688
rect 1273 712 1307 1688
rect 1431 712 1465 1688
rect 1689 712 1723 1688
rect -1611 619 -1543 653
rect -1396 619 -1342 653
rect -1195 619 -1127 653
rect -937 619 -869 653
rect -679 619 -611 653
rect -421 619 -353 653
rect -163 619 -95 653
rect 95 619 163 653
rect 353 619 421 653
rect 611 619 679 653
rect 869 619 937 653
rect 1127 619 1195 653
rect 1342 619 1396 653
rect 1543 619 1611 653
rect -1262 517 -1212 567
rect 1202 517 1252 567
rect 2822 423 2922 4117
rect -2822 118 -2760 218
rect -2760 118 2760 218
rect 2760 118 2822 218
rect -2822 -218 -2760 -118
rect -2760 -218 2760 -118
rect 2760 -218 2822 -118
rect -2922 -4117 -2822 -423
rect -41 -538 39 -458
rect -1611 -662 -1543 -628
rect -1396 -662 -1342 -628
rect -1195 -662 -1127 -628
rect -937 -662 -869 -628
rect -679 -662 -611 -628
rect -421 -662 -353 -628
rect -163 -662 -95 -628
rect 95 -662 163 -628
rect 353 -662 421 -628
rect 611 -662 679 -628
rect 869 -662 937 -628
rect 1127 -662 1195 -628
rect 1342 -662 1396 -628
rect 1543 -662 1611 -628
rect -1723 -1688 -1689 -712
rect -1465 -1688 -1431 -712
rect -1307 -1688 -1273 -712
rect -1049 -1688 -1015 -712
rect -791 -1688 -757 -712
rect -533 -1688 -499 -712
rect -275 -1688 -241 -712
rect -17 -1688 17 -712
rect 241 -1688 275 -712
rect 499 -1688 533 -712
rect 757 -1688 791 -712
rect 1015 -1688 1049 -712
rect 1273 -1688 1307 -712
rect 1431 -1688 1465 -712
rect 1689 -1688 1723 -712
rect -1611 -1772 -1543 -1738
rect -1396 -1772 -1342 -1738
rect -1195 -1772 -1127 -1738
rect -937 -1772 -869 -1738
rect -679 -1772 -611 -1738
rect -421 -1772 -353 -1738
rect -163 -1772 -95 -1738
rect 95 -1772 163 -1738
rect 353 -1772 421 -1738
rect 611 -1772 679 -1738
rect 869 -1772 937 -1738
rect 1127 -1772 1195 -1738
rect 1342 -1772 1396 -1738
rect 1543 -1772 1611 -1738
rect -685 -1902 -605 -1822
rect -427 -1902 -347 -1822
rect 347 -1902 427 -1822
rect 605 -1902 685 -1822
rect -556 -2126 -476 -2046
rect 476 -2126 556 -2046
rect -2227 -2462 -2159 -2428
rect -1969 -2462 -1901 -2428
rect -1711 -2462 -1643 -2428
rect -1453 -2462 -1385 -2428
rect -1195 -2462 -1127 -2428
rect -937 -2462 -869 -2428
rect -679 -2462 -611 -2428
rect -421 -2462 -353 -2428
rect -163 -2462 -95 -2428
rect 95 -2462 163 -2428
rect 353 -2462 421 -2428
rect 611 -2462 679 -2428
rect 869 -2462 937 -2428
rect 1127 -2462 1195 -2428
rect 1385 -2462 1453 -2428
rect 1643 -2462 1711 -2428
rect 1901 -2462 1969 -2428
rect 2159 -2462 2227 -2428
rect -2339 -3488 -2305 -2512
rect -2081 -3488 -2047 -2512
rect -1823 -3488 -1789 -2512
rect -1565 -3488 -1531 -2512
rect -1307 -3488 -1273 -2512
rect -1049 -3488 -1015 -2512
rect -791 -3488 -757 -2512
rect -533 -3488 -499 -2512
rect -275 -3488 -241 -2512
rect -17 -3488 17 -2512
rect 241 -3488 275 -2512
rect 499 -3488 533 -2512
rect 757 -3488 791 -2512
rect 1015 -3488 1049 -2512
rect 1273 -3488 1307 -2512
rect 1531 -3488 1565 -2512
rect 1789 -3488 1823 -2512
rect 2047 -3488 2081 -2512
rect 2305 -3488 2339 -2512
rect -2227 -3572 -2159 -3538
rect -1969 -3572 -1901 -3538
rect -1711 -3572 -1643 -3538
rect -1453 -3572 -1385 -3538
rect -1195 -3572 -1127 -3538
rect -937 -3572 -869 -3538
rect -679 -3572 -611 -3538
rect -421 -3572 -353 -3538
rect -163 -3572 -95 -3538
rect 95 -3572 163 -3538
rect 353 -3572 421 -3538
rect 611 -3572 679 -3538
rect 869 -3572 937 -3538
rect 1127 -3572 1195 -3538
rect 1385 -3572 1453 -3538
rect 1643 -3572 1711 -3538
rect 1901 -3572 1969 -3538
rect 2159 -3572 2227 -3538
rect 2822 -4117 2922 -423
rect -2822 -4422 -2760 -4322
rect -2760 -4422 2760 -4322
rect 2760 -4422 2822 -4322
<< metal1 >>
rect -2928 4422 2928 4428
rect -2928 4322 -2822 4422
rect 2822 4322 2928 4422
rect -2928 4316 2928 4322
rect -2928 4117 -2816 4316
rect -2928 423 -2922 4117
rect -2822 3746 -2816 4117
rect -2216 4016 -2206 4316
rect 2206 4016 2216 4316
rect 2816 4117 2928 4316
rect 2816 3746 2822 4117
rect -2822 3654 -235 3746
rect -2822 2038 -2816 3654
rect -2345 3587 -2299 3654
rect -2345 3581 -2147 3587
rect -2345 3547 -2227 3581
rect -2159 3547 -2147 3581
rect -2345 3541 -2147 3547
rect -1981 3581 -1889 3587
rect -1981 3547 -1969 3581
rect -1901 3547 -1889 3581
rect -1981 3541 -1889 3547
rect -2345 3488 -2299 3541
rect -2345 2512 -2339 3488
rect -2305 2512 -2299 3488
rect -2345 2500 -2299 2512
rect -2087 3488 -2041 3500
rect -2087 2512 -2081 3488
rect -2047 2512 -2041 3488
rect -2087 2459 -2041 2512
rect -1829 3488 -1783 3654
rect -1313 3587 -1267 3654
rect -1723 3581 -1631 3587
rect -1723 3547 -1711 3581
rect -1643 3547 -1631 3581
rect -1723 3541 -1631 3547
rect -1465 3581 -1373 3587
rect -1465 3547 -1453 3581
rect -1385 3547 -1373 3581
rect -1465 3541 -1373 3547
rect -1313 3581 -1115 3587
rect -1313 3547 -1195 3581
rect -1127 3547 -1115 3581
rect -1313 3541 -1115 3547
rect -949 3581 -857 3587
rect -949 3547 -937 3581
rect -869 3547 -857 3581
rect -949 3541 -857 3547
rect -1829 2512 -1823 3488
rect -1789 2512 -1783 3488
rect -1829 2500 -1783 2512
rect -1571 3488 -1525 3500
rect -1571 2512 -1565 3488
rect -1531 2512 -1525 3488
rect -2239 2453 -2147 2459
rect -2239 2419 -2227 2453
rect -2159 2419 -2147 2453
rect -2239 2413 -2147 2419
rect -2087 2453 -1889 2459
rect -2087 2419 -1969 2453
rect -1901 2419 -1889 2453
rect -2087 2367 -1889 2419
rect -1723 2453 -1631 2459
rect -1723 2419 -1711 2453
rect -1643 2419 -1631 2453
rect -1723 2413 -1631 2419
rect -2087 2162 -2041 2367
rect -1571 2254 -1525 2512
rect -1313 3488 -1267 3541
rect -1313 2512 -1307 3488
rect -1273 2512 -1267 3488
rect -1313 2500 -1267 2512
rect -1055 3488 -1009 3500
rect -1055 2512 -1049 3488
rect -1015 2512 -1009 3488
rect -1055 2459 -1009 2512
rect -797 3488 -751 3654
rect -691 3581 -599 3587
rect -691 3547 -679 3581
rect -611 3547 -599 3581
rect -691 3541 -599 3547
rect -433 3581 -341 3587
rect -433 3547 -421 3581
rect -353 3547 -341 3581
rect -433 3541 -341 3547
rect -797 2512 -791 3488
rect -757 2512 -751 3488
rect -797 2500 -751 2512
rect -539 3488 -493 3500
rect -539 2512 -533 3488
rect -499 2512 -493 3488
rect -1465 2453 -1373 2459
rect -1465 2419 -1453 2453
rect -1385 2419 -1373 2453
rect -1465 2413 -1373 2419
rect -1207 2453 -1115 2459
rect -1207 2419 -1195 2453
rect -1127 2419 -1115 2453
rect -1207 2413 -1115 2419
rect -1055 2453 -857 2459
rect -1055 2419 -937 2453
rect -869 2419 -857 2453
rect -1055 2367 -857 2419
rect -691 2453 -599 2459
rect -691 2419 -679 2453
rect -611 2419 -599 2453
rect -691 2413 -599 2419
rect -1571 2248 -1507 2254
rect -1571 2196 -1565 2248
rect -1513 2196 -1507 2248
rect -1571 2190 -1507 2196
rect -1055 2162 -1009 2367
rect -539 2346 -493 2512
rect -281 3488 -235 3654
rect 235 3654 2822 3746
rect -175 3581 -83 3587
rect -175 3547 -163 3581
rect -95 3547 -83 3581
rect -175 3541 -83 3547
rect 83 3581 175 3587
rect 83 3547 95 3581
rect 163 3547 175 3581
rect 83 3541 175 3547
rect -281 2512 -275 3488
rect -241 2512 -235 3488
rect -281 2500 -235 2512
rect -23 3488 23 3500
rect -23 2512 -17 3488
rect 17 2512 23 3488
rect -23 2459 23 2512
rect 235 3488 281 3654
rect 341 3581 433 3587
rect 341 3547 353 3581
rect 421 3547 433 3581
rect 341 3541 433 3547
rect 599 3581 691 3587
rect 599 3547 611 3581
rect 679 3547 691 3581
rect 599 3541 691 3547
rect 235 2512 241 3488
rect 275 2512 281 3488
rect 235 2500 281 2512
rect 493 3488 539 3500
rect 493 2512 499 3488
rect 533 2512 539 3488
rect -433 2453 -341 2459
rect -433 2419 -421 2453
rect -353 2419 -341 2453
rect -433 2413 -341 2419
rect -175 2453 175 2459
rect -175 2419 -163 2453
rect -95 2450 95 2453
rect -95 2419 -54 2450
rect -175 2389 -54 2419
rect 55 2419 95 2450
rect 163 2419 175 2453
rect 55 2389 175 2419
rect 341 2453 433 2459
rect 341 2419 353 2453
rect 421 2419 433 2453
rect 341 2413 433 2419
rect -175 2380 175 2389
rect 493 2346 539 2512
rect 751 3488 797 3654
rect 1267 3587 1313 3654
rect 857 3581 949 3587
rect 857 3547 869 3581
rect 937 3547 949 3581
rect 857 3541 949 3547
rect 1115 3581 1313 3587
rect 1115 3547 1127 3581
rect 1195 3547 1313 3581
rect 1115 3541 1313 3547
rect 1373 3581 1465 3587
rect 1373 3547 1385 3581
rect 1453 3547 1465 3581
rect 1373 3541 1465 3547
rect 1631 3581 1723 3587
rect 1631 3547 1643 3581
rect 1711 3547 1723 3581
rect 1631 3541 1723 3547
rect 751 2512 757 3488
rect 791 2512 797 3488
rect 751 2500 797 2512
rect 1009 3488 1055 3500
rect 1009 2512 1015 3488
rect 1049 2512 1055 3488
rect 1009 2459 1055 2512
rect 1267 3488 1313 3541
rect 1267 2512 1273 3488
rect 1307 2512 1313 3488
rect 1267 2500 1313 2512
rect 1525 3488 1571 3500
rect 1525 2512 1531 3488
rect 1565 2512 1571 3488
rect 599 2453 691 2459
rect 599 2419 611 2453
rect 679 2419 691 2453
rect 599 2413 691 2419
rect 857 2453 1055 2459
rect 857 2419 869 2453
rect 937 2419 1055 2453
rect 857 2367 1055 2419
rect 1115 2453 1207 2459
rect 1115 2419 1127 2453
rect 1195 2419 1207 2453
rect 1115 2413 1207 2419
rect 1373 2453 1465 2459
rect 1373 2419 1385 2453
rect 1453 2419 1465 2453
rect 1373 2413 1465 2419
rect -539 2340 -475 2346
rect -671 2288 -567 2294
rect -671 2196 -665 2288
rect -573 2196 -567 2288
rect -539 2288 -533 2340
rect -481 2288 -475 2340
rect -539 2282 -475 2288
rect -33 2340 31 2346
rect -33 2288 -27 2340
rect 25 2288 31 2340
rect -671 2190 -567 2196
rect -2087 2156 -2023 2162
rect -2087 2104 -2081 2156
rect -2029 2104 -2023 2156
rect -2087 2098 -2023 2104
rect -1064 2156 -1000 2162
rect -1064 2104 -1058 2156
rect -1006 2104 -1000 2156
rect -1064 2098 -1000 2104
rect -2822 2010 -1115 2038
rect -2822 1890 -2816 2010
rect -2556 1976 -1238 1982
rect -2556 1924 -2550 1976
rect -2498 1924 -1238 1976
rect -2556 1918 -1238 1924
rect -1302 1912 -1238 1918
rect -2822 1826 -1436 1890
rect -2822 423 -2816 1826
rect -1471 1787 -1436 1826
rect -1302 1860 -1296 1912
rect -1244 1860 -1238 1912
rect -1302 1854 -1238 1860
rect -1729 1781 -1436 1787
rect -1729 1747 -1611 1781
rect -1543 1747 -1436 1781
rect -1729 1741 -1436 1747
rect -1408 1781 -1330 1787
rect -1408 1747 -1396 1781
rect -1342 1747 -1330 1781
rect -1408 1741 -1330 1747
rect -1729 1688 -1683 1741
rect -1729 712 -1723 1688
rect -1689 712 -1683 1688
rect -1729 700 -1683 712
rect -1471 1700 -1436 1741
rect -1302 1700 -1267 1854
rect -1207 1781 -1115 2010
rect -975 2014 -901 2020
rect -975 1952 -969 2014
rect -907 1952 -901 2014
rect -975 1946 -901 1952
rect -797 2004 -733 2010
rect -797 1952 -791 2004
rect -739 1952 -733 2004
rect -797 1946 -733 1952
rect -290 2003 -226 2009
rect -290 1951 -284 2003
rect -232 1951 -226 2003
rect -1207 1747 -1195 1781
rect -1127 1747 -1115 1781
rect -1207 1741 -1115 1747
rect -949 1781 -857 1787
rect -949 1747 -937 1781
rect -869 1747 -857 1781
rect -949 1741 -857 1747
rect -1471 1688 -1425 1700
rect -1471 712 -1465 1688
rect -1431 712 -1425 1688
rect -1471 700 -1425 712
rect -1313 1688 -1267 1700
rect -1313 712 -1307 1688
rect -1273 712 -1267 1688
rect -1313 700 -1267 712
rect -1055 1688 -1009 1700
rect -1055 712 -1049 1688
rect -1015 712 -1009 1688
rect -1623 653 -1531 659
rect -1623 619 -1611 653
rect -1543 619 -1531 653
rect -1623 613 -1531 619
rect -1408 653 -1330 659
rect -1408 619 -1396 653
rect -1342 619 -1330 653
rect -1408 613 -1330 619
rect -1207 653 -1115 659
rect -1207 619 -1195 653
rect -1127 619 -1115 653
rect -1207 613 -1115 619
rect -1274 573 -1200 579
rect -1274 511 -1268 573
rect -1206 511 -1200 573
rect -1274 505 -1200 511
rect -1055 546 -1009 712
rect -797 1688 -751 1946
rect -290 1945 -226 1951
rect -33 2004 31 2288
rect 475 2340 539 2346
rect 475 2288 481 2340
rect 533 2288 539 2340
rect 475 2282 539 2288
rect 567 2288 671 2294
rect 567 2196 573 2288
rect 665 2196 671 2288
rect 567 2190 671 2196
rect 1009 2162 1055 2367
rect 1525 2254 1571 2512
rect 1783 3488 1829 3654
rect 2299 3587 2345 3654
rect 1889 3581 1981 3587
rect 1889 3547 1901 3581
rect 1969 3547 1981 3581
rect 1889 3541 1981 3547
rect 2147 3581 2345 3587
rect 2147 3547 2159 3581
rect 2227 3547 2345 3581
rect 2147 3541 2345 3547
rect 1783 2512 1789 3488
rect 1823 2512 1829 3488
rect 1783 2500 1829 2512
rect 2041 3488 2087 3500
rect 2041 2512 2047 3488
rect 2081 2512 2087 3488
rect 2041 2459 2087 2512
rect 2299 3488 2345 3541
rect 2299 2512 2305 3488
rect 2339 2512 2345 3488
rect 2299 2500 2345 2512
rect 1631 2453 1723 2459
rect 1631 2419 1643 2453
rect 1711 2419 1723 2453
rect 1631 2413 1723 2419
rect 1889 2453 2087 2459
rect 1889 2419 1901 2453
rect 1969 2419 2087 2453
rect 1889 2367 2087 2419
rect 2147 2453 2239 2459
rect 2147 2419 2159 2453
rect 2227 2419 2239 2453
rect 2147 2413 2239 2419
rect 1507 2248 1571 2254
rect 1507 2196 1513 2248
rect 1565 2196 1571 2248
rect 1507 2190 1571 2196
rect 2041 2162 2087 2367
rect 1000 2156 1064 2162
rect 1000 2104 1006 2156
rect 1058 2104 1064 2156
rect 1000 2098 1064 2104
rect 2023 2156 2087 2162
rect 2023 2104 2029 2156
rect 2081 2104 2087 2156
rect 2023 2098 2087 2104
rect 2816 2038 2822 3654
rect 901 2014 975 2020
rect -33 1952 -27 2004
rect 25 1952 31 2004
rect -33 1945 31 1952
rect 226 2004 290 2010
rect 226 1952 232 2004
rect 284 1952 290 2004
rect 226 1946 290 1952
rect 733 2004 797 2010
rect 733 1952 739 2004
rect 791 1952 797 2004
rect 733 1946 797 1952
rect 901 1952 907 2014
rect 969 1952 975 2014
rect 901 1946 975 1952
rect 1115 2010 2822 2038
rect -691 1781 -599 1787
rect -691 1747 -679 1781
rect -611 1747 -599 1781
rect -691 1741 -599 1747
rect -433 1781 -341 1787
rect -433 1747 -421 1781
rect -353 1747 -341 1781
rect -433 1741 -341 1747
rect -797 712 -791 1688
rect -757 712 -751 1688
rect -797 700 -751 712
rect -539 1688 -493 1700
rect -539 712 -533 1688
rect -499 712 -493 1688
rect -949 653 -857 659
rect -949 619 -937 653
rect -869 619 -857 653
rect -949 613 -857 619
rect -691 653 -599 659
rect -691 619 -679 653
rect -611 619 -599 653
rect -691 613 -599 619
rect -1055 540 -991 546
rect -1055 488 -1049 540
rect -997 488 -991 540
rect -1055 482 -991 488
rect -2928 224 -2816 423
rect -539 362 -493 712
rect -281 1688 -235 1945
rect -175 1781 -83 1787
rect -175 1747 -163 1781
rect -95 1747 -83 1781
rect -175 1741 -83 1747
rect 83 1781 175 1787
rect 83 1747 95 1781
rect 163 1747 175 1781
rect 83 1741 175 1747
rect -281 712 -275 1688
rect -241 712 -235 1688
rect -281 700 -235 712
rect -23 1688 23 1700
rect -23 712 -17 1688
rect 17 712 23 1688
rect -433 653 -341 659
rect -433 619 -421 653
rect -353 619 -341 653
rect -433 613 -341 619
rect -175 653 -83 659
rect -175 619 -163 653
rect -95 619 -83 653
rect -175 613 -83 619
rect -23 546 23 712
rect 235 1688 281 1946
rect 341 1781 433 1787
rect 341 1747 353 1781
rect 421 1747 433 1781
rect 341 1741 433 1747
rect 599 1781 691 1787
rect 599 1747 611 1781
rect 679 1747 691 1781
rect 599 1741 691 1747
rect 235 712 241 1688
rect 275 712 281 1688
rect 235 700 281 712
rect 493 1688 539 1700
rect 493 712 499 1688
rect 533 712 539 1688
rect 83 653 175 659
rect 83 619 95 653
rect 163 619 175 653
rect 83 613 175 619
rect 341 653 433 659
rect 341 619 353 653
rect 421 619 433 653
rect 341 613 433 619
rect -32 540 32 546
rect -32 488 -26 540
rect 26 488 32 540
rect -32 482 32 488
rect 493 362 539 712
rect 751 1688 797 1946
rect 857 1781 949 1787
rect 857 1747 869 1781
rect 937 1747 949 1781
rect 857 1741 949 1747
rect 1115 1781 1207 2010
rect 1238 1976 2551 1982
rect 1238 1924 2493 1976
rect 2545 1924 2551 1976
rect 1238 1918 2551 1924
rect 1238 1912 1302 1918
rect 1238 1860 1244 1912
rect 1296 1860 1302 1912
rect 2816 1890 2822 2010
rect 1238 1854 1302 1860
rect 1115 1747 1127 1781
rect 1195 1747 1207 1781
rect 1115 1741 1207 1747
rect 1267 1700 1302 1854
rect 1436 1826 2822 1890
rect 1436 1787 1471 1826
rect 1330 1781 1408 1787
rect 1330 1747 1342 1781
rect 1396 1747 1408 1781
rect 1330 1741 1408 1747
rect 1436 1781 1729 1787
rect 1436 1747 1543 1781
rect 1611 1747 1729 1781
rect 1436 1741 1729 1747
rect 1436 1700 1471 1741
rect 751 712 757 1688
rect 791 712 797 1688
rect 751 700 797 712
rect 1009 1688 1055 1700
rect 1009 712 1015 1688
rect 1049 712 1055 1688
rect 599 653 691 659
rect 599 619 611 653
rect 679 619 691 653
rect 599 613 691 619
rect 857 653 949 659
rect 857 619 869 653
rect 937 619 949 653
rect 857 613 949 619
rect 1009 546 1055 712
rect 1267 1688 1313 1700
rect 1267 712 1273 1688
rect 1307 712 1313 1688
rect 1267 700 1313 712
rect 1425 1688 1471 1700
rect 1425 712 1431 1688
rect 1465 712 1471 1688
rect 1425 700 1471 712
rect 1683 1688 1729 1741
rect 1683 712 1689 1688
rect 1723 712 1729 1688
rect 1683 700 1729 712
rect 1115 653 1207 659
rect 1115 619 1127 653
rect 1195 619 1207 653
rect 1115 613 1207 619
rect 1330 653 1408 659
rect 1330 619 1342 653
rect 1396 619 1408 653
rect 1330 613 1408 619
rect 1531 653 1623 659
rect 1531 619 1543 653
rect 1611 619 1623 653
rect 1531 613 1623 619
rect 991 540 1055 546
rect 991 488 997 540
rect 1049 488 1055 540
rect 1190 573 1264 579
rect 1190 511 1196 573
rect 1258 511 1264 573
rect 1190 505 1264 511
rect 991 482 1055 488
rect 2816 423 2822 1826
rect 2922 423 2928 4117
rect -2392 356 -475 362
rect -2392 304 -2386 356
rect -2334 304 -533 356
rect -481 304 -475 356
rect -2392 298 -475 304
rect 475 356 2391 362
rect 475 304 481 356
rect 533 304 2333 356
rect 2385 304 2391 356
rect 475 298 2391 304
rect 2816 224 2928 423
rect -2928 218 2928 224
rect -2928 118 -2822 218
rect 2822 118 2928 218
rect -2928 112 2928 118
rect -2928 -118 2928 -112
rect -2928 -218 -2822 -118
rect 2822 -218 2928 -118
rect -2928 -224 2928 -218
rect -2928 -252 -2816 -224
rect 2816 -252 2928 -224
rect -2928 -316 2928 -252
rect -2928 -423 -2816 -316
rect -2556 -360 -1672 -354
rect -2556 -412 -2550 -360
rect -2498 -412 -1730 -360
rect -1678 -412 -1672 -360
rect -2556 -418 -1672 -412
rect -2928 -4117 -2922 -423
rect -2822 -2166 -2816 -423
rect -1471 -622 -1436 -316
rect -1302 -360 -1238 -354
rect -1302 -412 -1296 -360
rect -1244 -412 -1238 -360
rect -1302 -418 -1238 -412
rect -1729 -628 -1436 -622
rect -1729 -662 -1611 -628
rect -1543 -662 -1436 -628
rect -1729 -668 -1436 -662
rect -1408 -628 -1330 -622
rect -1408 -662 -1396 -628
rect -1342 -662 -1330 -628
rect -1408 -668 -1330 -662
rect -1729 -712 -1683 -668
rect -1729 -1688 -1723 -712
rect -1689 -1688 -1683 -712
rect -1729 -1700 -1683 -1688
rect -1471 -700 -1436 -668
rect -1302 -700 -1267 -418
rect -1207 -628 -1115 -316
rect -1207 -662 -1195 -628
rect -1127 -662 -1115 -628
rect -1207 -668 -1115 -662
rect -949 -628 -857 -622
rect -949 -662 -937 -628
rect -869 -662 -857 -628
rect -949 -668 -857 -662
rect -1471 -712 -1425 -700
rect -1471 -1688 -1465 -712
rect -1431 -1688 -1425 -712
rect -1471 -1700 -1425 -1688
rect -1313 -712 -1267 -700
rect -1313 -1688 -1307 -712
rect -1273 -1688 -1267 -712
rect -1313 -1700 -1267 -1688
rect -1055 -712 -1009 -700
rect -1055 -1688 -1049 -712
rect -1015 -1688 -1009 -712
rect -1623 -1738 -1531 -1732
rect -1623 -1772 -1611 -1738
rect -1543 -1772 -1531 -1738
rect -1623 -1778 -1531 -1772
rect -1408 -1738 -1330 -1732
rect -1408 -1772 -1396 -1738
rect -1342 -1772 -1330 -1738
rect -1408 -1778 -1330 -1772
rect -1207 -1738 -1115 -1732
rect -1207 -1772 -1195 -1738
rect -1127 -1772 -1115 -1738
rect -1207 -1778 -1115 -1772
rect -2556 -1856 -1836 -1850
rect -2556 -1908 -2550 -1856
rect -2498 -1908 -1894 -1856
rect -1842 -1908 -1836 -1856
rect -2556 -1914 -1836 -1908
rect -1055 -2034 -1009 -1688
rect -797 -712 -751 -316
rect -691 -628 -599 -622
rect -691 -662 -679 -628
rect -611 -662 -599 -628
rect -691 -668 -599 -662
rect -433 -628 -341 -622
rect -433 -662 -421 -628
rect -353 -662 -341 -628
rect -433 -668 -341 -662
rect -797 -1688 -791 -712
rect -757 -1688 -751 -712
rect -797 -1700 -751 -1688
rect -539 -712 -493 -700
rect -539 -1688 -533 -712
rect -499 -1688 -493 -712
rect -949 -1738 -857 -1732
rect -949 -1772 -937 -1738
rect -869 -1772 -857 -1738
rect -949 -1778 -857 -1772
rect -691 -1738 -599 -1732
rect -691 -1772 -679 -1738
rect -611 -1772 -599 -1738
rect -691 -1778 -599 -1772
rect -697 -1816 -593 -1810
rect -697 -1908 -691 -1816
rect -599 -1908 -593 -1816
rect -697 -1914 -593 -1908
rect -539 -1942 -493 -1688
rect -281 -712 -235 -316
rect -199 -360 207 -354
rect -199 -412 -193 -360
rect -141 -412 149 -360
rect 201 -412 207 -360
rect -199 -418 207 -412
rect -53 -452 51 -446
rect -53 -544 -47 -452
rect 45 -544 51 -452
rect -53 -550 51 -544
rect -175 -628 -83 -622
rect -175 -662 -163 -628
rect -95 -662 -83 -628
rect -175 -668 -83 -662
rect 83 -628 175 -622
rect 83 -662 95 -628
rect 163 -662 175 -628
rect 83 -668 175 -662
rect -281 -1688 -275 -712
rect -241 -1688 -235 -712
rect -281 -1700 -235 -1688
rect -23 -712 23 -700
rect -23 -1688 -17 -712
rect 17 -1688 23 -712
rect -433 -1738 -341 -1732
rect -433 -1772 -421 -1738
rect -353 -1772 -341 -1738
rect -433 -1778 -341 -1772
rect -175 -1738 -83 -1732
rect -175 -1772 -163 -1738
rect -95 -1772 -83 -1738
rect -175 -1778 -83 -1772
rect -439 -1816 -335 -1810
rect -439 -1908 -433 -1816
rect -341 -1908 -335 -1816
rect -439 -1914 -335 -1908
rect -539 -1948 -475 -1942
rect -539 -2000 -533 -1948
rect -481 -2000 -475 -1948
rect -539 -2006 -475 -2000
rect -23 -2034 23 -1688
rect 235 -712 281 -316
rect 341 -628 433 -622
rect 341 -662 353 -628
rect 421 -662 433 -628
rect 341 -668 433 -662
rect 599 -628 691 -622
rect 599 -662 611 -628
rect 679 -662 691 -628
rect 599 -668 691 -662
rect 235 -1688 241 -712
rect 275 -1688 281 -712
rect 235 -1700 281 -1688
rect 493 -712 539 -700
rect 493 -1688 499 -712
rect 533 -1688 539 -712
rect 83 -1738 175 -1732
rect 83 -1772 95 -1738
rect 163 -1772 175 -1738
rect 83 -1778 175 -1772
rect 341 -1738 433 -1732
rect 341 -1772 353 -1738
rect 421 -1772 433 -1738
rect 341 -1778 433 -1772
rect 335 -1816 439 -1810
rect 335 -1908 341 -1816
rect 433 -1908 439 -1816
rect 335 -1914 439 -1908
rect 493 -1942 539 -1688
rect 751 -712 797 -316
rect 857 -628 949 -622
rect 857 -662 869 -628
rect 937 -662 949 -628
rect 857 -668 949 -662
rect 1115 -628 1207 -316
rect 1238 -360 1302 -354
rect 1238 -412 1244 -360
rect 1296 -412 1302 -360
rect 1238 -418 1302 -412
rect 1115 -662 1127 -628
rect 1195 -662 1207 -628
rect 1115 -668 1207 -662
rect 1267 -700 1302 -418
rect 1436 -622 1471 -316
rect 1671 -360 2551 -354
rect 1671 -412 1677 -360
rect 1729 -412 2493 -360
rect 2545 -412 2551 -360
rect 1671 -418 2551 -412
rect 2816 -423 2928 -316
rect 1330 -628 1408 -622
rect 1330 -662 1342 -628
rect 1396 -662 1408 -628
rect 1330 -668 1408 -662
rect 1436 -628 1729 -622
rect 1436 -662 1543 -628
rect 1611 -662 1729 -628
rect 1436 -668 1729 -662
rect 1436 -700 1471 -668
rect 751 -1688 757 -712
rect 791 -1688 797 -712
rect 751 -1700 797 -1688
rect 1009 -712 1055 -700
rect 1009 -1688 1015 -712
rect 1049 -1688 1055 -712
rect 599 -1738 691 -1732
rect 599 -1772 611 -1738
rect 679 -1772 691 -1738
rect 599 -1778 691 -1772
rect 857 -1738 949 -1732
rect 857 -1772 869 -1738
rect 937 -1772 949 -1738
rect 857 -1778 949 -1772
rect 593 -1816 697 -1810
rect 593 -1908 599 -1816
rect 691 -1908 697 -1816
rect 593 -1914 697 -1908
rect 475 -1948 539 -1942
rect 475 -2000 481 -1948
rect 533 -2000 539 -1948
rect 475 -2006 539 -2000
rect 1009 -2034 1055 -1688
rect 1267 -712 1313 -700
rect 1267 -1688 1273 -712
rect 1307 -1688 1313 -712
rect 1267 -1700 1313 -1688
rect 1425 -712 1471 -700
rect 1425 -1688 1431 -712
rect 1465 -1688 1471 -712
rect 1425 -1700 1471 -1688
rect 1683 -712 1729 -668
rect 1683 -1688 1689 -712
rect 1723 -1688 1729 -712
rect 1683 -1700 1729 -1688
rect 1115 -1738 1207 -1732
rect 1115 -1772 1127 -1738
rect 1195 -1772 1207 -1738
rect 1115 -1778 1207 -1772
rect 1330 -1738 1408 -1732
rect 1330 -1772 1342 -1738
rect 1396 -1772 1408 -1738
rect 1330 -1778 1408 -1772
rect 1531 -1738 1623 -1732
rect 1531 -1772 1543 -1738
rect 1611 -1772 1623 -1738
rect 1531 -1778 1623 -1772
rect 1835 -1856 2555 -1850
rect 1835 -1908 1841 -1856
rect 1893 -1908 2497 -1856
rect 2549 -1908 2555 -1856
rect 1835 -1914 2555 -1908
rect -1055 -2040 -991 -2034
rect -1055 -2092 -1049 -2040
rect -997 -2092 -991 -2040
rect -1055 -2098 -991 -2092
rect -568 -2040 -464 -2034
rect -568 -2132 -562 -2040
rect -470 -2132 -464 -2040
rect -32 -2040 32 -2034
rect -32 -2092 -26 -2040
rect 26 -2092 32 -2040
rect -32 -2098 32 -2092
rect 464 -2040 568 -2034
rect -568 -2138 -464 -2132
rect 464 -2132 470 -2040
rect 562 -2132 568 -2040
rect 991 -2040 1055 -2034
rect 991 -2092 997 -2040
rect 1049 -2092 1055 -2040
rect 991 -2098 1055 -2092
rect 464 -2138 568 -2132
rect 2816 -2166 2822 -423
rect -2822 -2230 2822 -2166
rect -2822 -4117 -2816 -2230
rect -2239 -2428 -2147 -2230
rect -2096 -2316 -2032 -2310
rect -2096 -2368 -2090 -2316
rect -2038 -2368 -2032 -2316
rect -2096 -2374 -2032 -2368
rect -2345 -2462 -2227 -2428
rect -2159 -2462 -2147 -2428
rect -2345 -2468 -2147 -2462
rect -2345 -2512 -2299 -2468
rect -2345 -3488 -2339 -2512
rect -2305 -3488 -2299 -2512
rect -2345 -3500 -2299 -3488
rect -2087 -2512 -2041 -2374
rect -1981 -2428 -1889 -2422
rect -1981 -2462 -1969 -2428
rect -1901 -2462 -1889 -2428
rect -1981 -2468 -1889 -2462
rect -2087 -3488 -2081 -2512
rect -2047 -3488 -2041 -2512
rect -2087 -3500 -2041 -3488
rect -1829 -2512 -1783 -2230
rect -1723 -2316 -1631 -2310
rect -1723 -2368 -1717 -2316
rect -1637 -2368 -1631 -2316
rect -1723 -2428 -1631 -2368
rect -1723 -2462 -1711 -2428
rect -1643 -2462 -1631 -2428
rect -1723 -2468 -1631 -2462
rect -1465 -2316 -1373 -2310
rect -1465 -2368 -1459 -2316
rect -1379 -2368 -1373 -2316
rect -1465 -2428 -1373 -2368
rect -1465 -2462 -1453 -2428
rect -1385 -2462 -1373 -2428
rect -1465 -2468 -1373 -2462
rect -1829 -3488 -1823 -2512
rect -1789 -3488 -1783 -2512
rect -1829 -3500 -1783 -3488
rect -1571 -2512 -1525 -2500
rect -1571 -3488 -1565 -2512
rect -1531 -3488 -1525 -2512
rect -2239 -3538 -2147 -3532
rect -2239 -3572 -2227 -3538
rect -2159 -3572 -2147 -3538
rect -2239 -3578 -2147 -3572
rect -1981 -3538 -1889 -3532
rect -1981 -3572 -1969 -3538
rect -1901 -3572 -1889 -3538
rect -1981 -3632 -1889 -3572
rect -1723 -3538 -1631 -3532
rect -1723 -3572 -1711 -3538
rect -1643 -3572 -1631 -3538
rect -1723 -3578 -1631 -3572
rect -1571 -3626 -1525 -3488
rect -1313 -2512 -1267 -2230
rect -1064 -2316 -1000 -2310
rect -1064 -2368 -1058 -2316
rect -1006 -2368 -1000 -2316
rect -1064 -2374 -1000 -2368
rect -1207 -2428 -1115 -2422
rect -1207 -2462 -1195 -2428
rect -1127 -2462 -1115 -2428
rect -1207 -2468 -1115 -2462
rect -1313 -3488 -1307 -2512
rect -1273 -3488 -1267 -2512
rect -1313 -3500 -1267 -3488
rect -1055 -2512 -1009 -2374
rect -949 -2428 -857 -2230
rect -949 -2462 -937 -2428
rect -869 -2462 -857 -2428
rect -949 -2468 -857 -2462
rect -691 -2428 -599 -2422
rect -691 -2462 -679 -2428
rect -611 -2462 -599 -2428
rect -691 -2468 -599 -2462
rect -1055 -3488 -1049 -2512
rect -1015 -3488 -1009 -2512
rect -1055 -3500 -1009 -3488
rect -797 -2512 -751 -2500
rect -797 -3488 -791 -2512
rect -757 -3488 -751 -2512
rect -797 -3532 -751 -3488
rect -539 -2512 -493 -2230
rect -433 -2316 -341 -2310
rect -433 -2368 -427 -2316
rect -347 -2368 -341 -2316
rect -433 -2412 -341 -2368
rect -290 -2316 -226 -2310
rect -290 -2368 -284 -2316
rect -232 -2368 -226 -2316
rect -290 -2374 -226 -2368
rect -175 -2316 -83 -2310
rect -175 -2368 -169 -2316
rect -89 -2368 -83 -2316
rect -281 -2412 -235 -2374
rect -175 -2412 -83 -2368
rect -433 -2428 -83 -2412
rect -433 -2462 -421 -2428
rect -353 -2462 -163 -2428
rect -95 -2462 -83 -2428
rect -433 -2468 -83 -2462
rect -539 -3488 -533 -2512
rect -499 -3488 -493 -2512
rect -539 -3500 -493 -3488
rect -281 -2512 -235 -2468
rect -281 -3488 -275 -2512
rect -241 -3488 -235 -2512
rect -281 -3500 -235 -3488
rect -23 -2512 23 -2230
rect 83 -2428 175 -2422
rect 83 -2462 95 -2428
rect 163 -2462 175 -2428
rect 83 -2468 175 -2462
rect 341 -2428 433 -2422
rect 341 -2462 353 -2428
rect 421 -2462 433 -2428
rect 341 -2468 433 -2462
rect -23 -3488 -17 -2512
rect 17 -3488 23 -2512
rect -23 -3500 23 -3488
rect 235 -2512 281 -2500
rect 235 -3488 241 -2512
rect 275 -3488 281 -2512
rect 235 -3532 281 -3488
rect 493 -2512 539 -2230
rect 599 -2316 691 -2310
rect 599 -2368 605 -2316
rect 685 -2368 691 -2316
rect 599 -2412 691 -2368
rect 742 -2316 806 -2310
rect 742 -2368 748 -2316
rect 800 -2368 806 -2316
rect 742 -2374 806 -2368
rect 751 -2412 797 -2374
rect 599 -2428 797 -2412
rect 599 -2462 611 -2428
rect 679 -2462 797 -2428
rect 599 -2468 797 -2462
rect 857 -2428 949 -2230
rect 1000 -2316 1064 -2310
rect 1000 -2368 1006 -2316
rect 1058 -2368 1064 -2316
rect 1000 -2374 1064 -2368
rect 857 -2462 869 -2428
rect 937 -2462 949 -2428
rect 857 -2468 949 -2462
rect 493 -3488 499 -2512
rect 533 -3488 539 -2512
rect 493 -3500 539 -3488
rect 751 -2512 797 -2468
rect 751 -3488 757 -2512
rect 791 -3488 797 -2512
rect 751 -3500 797 -3488
rect 1009 -2512 1055 -2374
rect 1115 -2428 1207 -2422
rect 1115 -2462 1127 -2428
rect 1195 -2462 1207 -2428
rect 1115 -2468 1207 -2462
rect 1009 -3488 1015 -2512
rect 1049 -3488 1055 -2512
rect 1009 -3500 1055 -3488
rect 1267 -2512 1313 -2230
rect 1373 -2316 1465 -2310
rect 1373 -2368 1379 -2316
rect 1459 -2368 1465 -2316
rect 1373 -2428 1465 -2368
rect 1373 -2462 1385 -2428
rect 1453 -2462 1465 -2428
rect 1373 -2468 1465 -2462
rect 1631 -2316 1723 -2310
rect 1631 -2368 1637 -2316
rect 1717 -2368 1723 -2316
rect 1631 -2428 1723 -2368
rect 1631 -2462 1643 -2428
rect 1711 -2462 1723 -2428
rect 1631 -2468 1723 -2462
rect 1267 -3488 1273 -2512
rect 1307 -3488 1313 -2512
rect 1267 -3500 1313 -3488
rect 1525 -2512 1571 -2500
rect 1525 -3488 1531 -2512
rect 1565 -3488 1571 -2512
rect -1465 -3538 -1373 -3532
rect -1465 -3572 -1453 -3538
rect -1385 -3572 -1373 -3538
rect -1465 -3578 -1373 -3572
rect -1207 -3538 -1115 -3532
rect -1207 -3572 -1195 -3538
rect -1127 -3572 -1115 -3538
rect -1981 -3684 -1975 -3632
rect -1895 -3684 -1889 -3632
rect -1981 -3690 -1889 -3684
rect -1580 -3632 -1516 -3626
rect -1580 -3684 -1574 -3632
rect -1522 -3684 -1516 -3632
rect -1580 -3690 -1516 -3684
rect -1207 -3632 -1115 -3572
rect -949 -3538 -857 -3532
rect -949 -3572 -937 -3538
rect -869 -3572 -857 -3538
rect -949 -3578 -857 -3572
rect -797 -3538 -599 -3532
rect -797 -3572 -679 -3538
rect -611 -3572 -599 -3538
rect -797 -3588 -599 -3572
rect -433 -3538 -341 -3532
rect -433 -3572 -421 -3538
rect -353 -3572 -341 -3538
rect -433 -3578 -341 -3572
rect -175 -3538 -83 -3532
rect -175 -3572 -163 -3538
rect -95 -3572 -83 -3538
rect -175 -3578 -83 -3572
rect 83 -3538 433 -3532
rect 83 -3572 95 -3538
rect 163 -3572 353 -3538
rect 421 -3572 433 -3538
rect -797 -3626 -751 -3588
rect -1207 -3684 -1201 -3632
rect -1121 -3684 -1115 -3632
rect -1207 -3690 -1115 -3684
rect -806 -3632 -742 -3626
rect -806 -3684 -800 -3632
rect -748 -3684 -742 -3632
rect -806 -3690 -742 -3684
rect -691 -3632 -599 -3588
rect -691 -3684 -685 -3632
rect -605 -3684 -599 -3632
rect -691 -3690 -599 -3684
rect 83 -3589 433 -3572
rect 599 -3538 691 -3532
rect 599 -3572 611 -3538
rect 679 -3572 691 -3538
rect 599 -3578 691 -3572
rect 857 -3538 949 -3532
rect 857 -3572 869 -3538
rect 937 -3572 949 -3538
rect 857 -3578 949 -3572
rect 1115 -3538 1207 -3532
rect 1115 -3572 1127 -3538
rect 1195 -3572 1207 -3538
rect 83 -3632 175 -3589
rect 235 -3626 281 -3589
rect 83 -3684 89 -3632
rect 169 -3684 175 -3632
rect 83 -3690 175 -3684
rect 226 -3632 290 -3626
rect 226 -3684 232 -3632
rect 284 -3684 290 -3632
rect 226 -3690 290 -3684
rect 341 -3632 433 -3589
rect 341 -3684 347 -3632
rect 427 -3684 433 -3632
rect 341 -3690 433 -3684
rect 1115 -3632 1207 -3572
rect 1373 -3538 1465 -3532
rect 1373 -3572 1385 -3538
rect 1453 -3572 1465 -3538
rect 1373 -3578 1465 -3572
rect 1525 -3626 1571 -3488
rect 1783 -2512 1829 -2230
rect 2032 -2316 2096 -2310
rect 2032 -2368 2038 -2316
rect 2090 -2368 2096 -2316
rect 2032 -2374 2096 -2368
rect 1889 -2428 1981 -2422
rect 1889 -2462 1901 -2428
rect 1969 -2462 1981 -2428
rect 1889 -2468 1981 -2462
rect 1783 -3488 1789 -2512
rect 1823 -3488 1829 -2512
rect 1783 -3500 1829 -3488
rect 2041 -2512 2087 -2374
rect 2147 -2428 2239 -2230
rect 2147 -2462 2159 -2428
rect 2227 -2462 2345 -2428
rect 2147 -2468 2345 -2462
rect 2041 -3488 2047 -2512
rect 2081 -3488 2087 -2512
rect 2041 -3500 2087 -3488
rect 2299 -2512 2345 -2468
rect 2299 -3488 2305 -2512
rect 2339 -3488 2345 -2512
rect 2299 -3500 2345 -3488
rect 1631 -3538 1723 -3532
rect 1631 -3572 1643 -3538
rect 1711 -3572 1723 -3538
rect 1631 -3578 1723 -3572
rect 1889 -3538 1981 -3532
rect 1889 -3572 1901 -3538
rect 1969 -3572 1981 -3538
rect 1115 -3684 1121 -3632
rect 1201 -3684 1207 -3632
rect 1115 -3690 1207 -3684
rect 1516 -3632 1580 -3626
rect 1516 -3684 1522 -3632
rect 1574 -3684 1580 -3632
rect 1516 -3690 1580 -3684
rect 1889 -3632 1981 -3572
rect 2147 -3538 2239 -3532
rect 2147 -3572 2159 -3538
rect 2227 -3572 2239 -3538
rect 2147 -3578 2239 -3572
rect 1889 -3684 1895 -3632
rect 1975 -3684 1981 -3632
rect 1889 -3690 1981 -3684
rect -2928 -4316 -2816 -4117
rect -2216 -4316 -2206 -4016
rect 2206 -4316 2216 -4016
rect 2816 -4117 2822 -2230
rect 2922 -4117 2928 -423
rect 2816 -4316 2928 -4117
rect -2928 -4322 2928 -4316
rect -2928 -4422 -2822 -4322
rect 2822 -4422 2928 -4322
rect -2928 -4428 2928 -4422
<< via1 >>
rect -2816 4016 -2216 4316
rect 2216 4016 2816 4316
rect -1565 2196 -1513 2248
rect -54 2389 55 2450
rect -665 2282 -573 2288
rect -665 2202 -659 2282
rect -659 2202 -579 2282
rect -579 2202 -573 2282
rect -665 2196 -573 2202
rect -533 2288 -481 2340
rect -27 2288 25 2340
rect -2081 2104 -2029 2156
rect -1058 2104 -1006 2156
rect -2550 1924 -2498 1976
rect -1296 1860 -1244 1912
rect -969 2008 -907 2014
rect -969 1958 -963 2008
rect -963 1958 -913 2008
rect -913 1958 -907 2008
rect -969 1952 -907 1958
rect -791 1952 -739 2004
rect -284 1951 -232 2003
rect -1268 567 -1206 573
rect -1268 517 -1262 567
rect -1262 517 -1212 567
rect -1212 517 -1206 567
rect -1268 511 -1206 517
rect 481 2288 533 2340
rect 573 2282 665 2288
rect 573 2202 579 2282
rect 579 2202 659 2282
rect 659 2202 665 2282
rect 573 2196 665 2202
rect 1513 2196 1565 2248
rect 1006 2104 1058 2156
rect 2029 2104 2081 2156
rect -27 1952 25 2004
rect 232 1952 284 2004
rect 739 1952 791 2004
rect 907 2008 969 2014
rect 907 1958 913 2008
rect 913 1958 963 2008
rect 963 1958 969 2008
rect 907 1952 969 1958
rect -1049 488 -997 540
rect -26 488 26 540
rect 2493 1924 2545 1976
rect 1244 1860 1296 1912
rect 997 488 1049 540
rect 1196 567 1258 573
rect 1196 517 1202 567
rect 1202 517 1252 567
rect 1252 517 1258 567
rect 1196 511 1258 517
rect -2386 304 -2334 356
rect -533 304 -481 356
rect 481 304 533 356
rect 2333 304 2385 356
rect -2550 -412 -2498 -360
rect -1730 -412 -1678 -360
rect -1296 -412 -1244 -360
rect -2550 -1908 -2498 -1856
rect -1894 -1908 -1842 -1856
rect -691 -1822 -599 -1816
rect -691 -1902 -685 -1822
rect -685 -1902 -605 -1822
rect -605 -1902 -599 -1822
rect -691 -1908 -599 -1902
rect -193 -412 -141 -360
rect 149 -412 201 -360
rect -47 -458 45 -452
rect -47 -538 -41 -458
rect -41 -538 39 -458
rect 39 -538 45 -458
rect -47 -544 45 -538
rect -433 -1822 -341 -1816
rect -433 -1902 -427 -1822
rect -427 -1902 -347 -1822
rect -347 -1902 -341 -1822
rect -433 -1908 -341 -1902
rect -533 -2000 -481 -1948
rect 341 -1822 433 -1816
rect 341 -1902 347 -1822
rect 347 -1902 427 -1822
rect 427 -1902 433 -1822
rect 341 -1908 433 -1902
rect 1244 -412 1296 -360
rect 1677 -412 1729 -360
rect 2493 -412 2545 -360
rect 599 -1822 691 -1816
rect 599 -1902 605 -1822
rect 605 -1902 685 -1822
rect 685 -1902 691 -1822
rect 599 -1908 691 -1902
rect 481 -2000 533 -1948
rect 1841 -1908 1893 -1856
rect 2497 -1908 2549 -1856
rect -1049 -2092 -997 -2040
rect -562 -2046 -470 -2040
rect -562 -2126 -556 -2046
rect -556 -2126 -476 -2046
rect -476 -2126 -470 -2046
rect -562 -2132 -470 -2126
rect -26 -2092 26 -2040
rect 470 -2046 562 -2040
rect 470 -2126 476 -2046
rect 476 -2126 556 -2046
rect 556 -2126 562 -2046
rect 470 -2132 562 -2126
rect 997 -2092 1049 -2040
rect -2090 -2368 -2038 -2316
rect -1717 -2368 -1637 -2316
rect -1459 -2368 -1379 -2316
rect -1058 -2368 -1006 -2316
rect -427 -2368 -347 -2316
rect -284 -2368 -232 -2316
rect -169 -2368 -89 -2316
rect 605 -2368 685 -2316
rect 748 -2368 800 -2316
rect 1006 -2368 1058 -2316
rect 1379 -2368 1459 -2316
rect 1637 -2368 1717 -2316
rect -1975 -3684 -1895 -3632
rect -1574 -3684 -1522 -3632
rect -1201 -3684 -1121 -3632
rect -800 -3684 -748 -3632
rect -685 -3684 -605 -3632
rect 89 -3684 169 -3632
rect 232 -3684 284 -3632
rect 347 -3684 427 -3632
rect 2038 -2368 2090 -2316
rect 1121 -3684 1201 -3632
rect 1522 -3684 1574 -3632
rect 1895 -3684 1975 -3632
rect -2816 -4316 -2216 -4016
rect 2216 -4316 2816 -4016
<< metal2 >>
rect -2816 4316 -2216 4326
rect -2816 4006 -2216 4016
rect 2216 4316 2816 4326
rect 2216 4006 2816 4016
rect -63 2450 63 2459
rect -63 2389 -54 2450
rect 55 2389 63 2450
rect -63 2380 63 2389
rect -539 2340 539 2346
rect -671 2288 -567 2294
rect -671 2254 -665 2288
rect -2228 2248 -665 2254
rect -2228 2196 -1565 2248
rect -1513 2196 -665 2248
rect -573 2254 -567 2288
rect -539 2288 -533 2340
rect -481 2288 -27 2340
rect 25 2288 481 2340
rect 533 2288 539 2340
rect -539 2282 539 2288
rect 567 2288 671 2294
rect 567 2254 573 2288
rect -573 2196 573 2254
rect 665 2254 671 2288
rect 665 2248 2227 2254
rect 665 2196 1513 2248
rect 1565 2196 2227 2248
rect -2228 2190 2227 2196
rect -2556 1976 -2492 1982
rect -2556 1924 -2550 1976
rect -2498 1924 -2492 1976
rect -2556 -360 -2492 1924
rect -2556 -412 -2550 -360
rect -2498 -412 -2492 -360
rect -2556 -418 -2492 -412
rect -2392 356 -2328 362
rect -2392 304 -2386 356
rect -2334 304 -2328 356
rect -2556 -1856 -2492 -1850
rect -2556 -1908 -2550 -1856
rect -2498 -1908 -2492 -1856
rect -2556 -3718 -2492 -1908
rect -2392 -2218 -2328 304
rect -2228 -2034 -2164 2190
rect -2087 2156 2087 2162
rect -2087 2104 -2081 2156
rect -2029 2104 -1058 2156
rect -1006 2104 1006 2156
rect 1058 2104 2029 2156
rect 2081 2104 2087 2156
rect -2087 2098 2087 2104
rect -1576 2070 -1512 2098
rect -2064 2006 -1512 2070
rect 1512 2070 1576 2098
rect -975 2014 -901 2020
rect -2064 -1942 -2000 2006
rect -975 1952 -969 2014
rect -907 1952 -901 2014
rect 901 2014 975 2020
rect -975 1946 -901 1952
rect -797 2004 797 2010
rect -797 1952 -791 2004
rect -739 2003 -27 2004
rect -739 1952 -284 2003
rect -797 1951 -284 1952
rect -232 1952 -27 2003
rect 25 1952 232 2004
rect 284 1952 739 2004
rect 791 1952 797 2004
rect -232 1951 797 1952
rect -797 1946 797 1951
rect 901 1952 907 2014
rect 969 1952 975 2014
rect 1512 2006 2063 2070
rect 901 1946 975 1952
rect -1302 1912 1302 1918
rect -1302 1860 -1296 1912
rect -1244 1860 1244 1912
rect 1296 1860 1302 1912
rect -1302 1854 1302 1860
rect -1274 573 -1200 579
rect -1274 511 -1268 573
rect -1206 511 -1200 573
rect 1190 573 1264 579
rect -1274 505 -1200 511
rect -1055 540 1055 546
rect -1055 488 -1049 540
rect -997 488 -26 540
rect 26 488 997 540
rect 1049 488 1055 540
rect 1190 511 1196 573
rect 1258 511 1264 573
rect 1190 505 1264 511
rect -1055 482 1055 488
rect -32 454 32 482
rect -1900 390 1899 454
rect -1900 -1850 -1836 390
rect -539 356 539 362
rect -539 304 -533 356
rect -481 304 481 356
rect 533 304 539 356
rect -539 298 539 304
rect -1736 -360 -135 -354
rect -1736 -412 -1730 -360
rect -1678 -412 -1296 -360
rect -1244 -412 -193 -360
rect -141 -412 -135 -360
rect -1736 -418 -135 -412
rect -33 -446 31 298
rect 143 -360 1735 -354
rect 143 -412 149 -360
rect 201 -412 1244 -360
rect 1296 -412 1677 -360
rect 1729 -412 1735 -360
rect 143 -418 1735 -412
rect -53 -452 51 -446
rect -53 -544 -47 -452
rect 45 -544 51 -452
rect -53 -550 51 -544
rect -697 -1816 -593 -1810
rect -697 -1850 -691 -1816
rect -1900 -1856 -691 -1850
rect -1900 -1908 -1894 -1856
rect -1842 -1908 -691 -1856
rect -599 -1850 -593 -1816
rect -439 -1816 -335 -1810
rect -439 -1850 -433 -1816
rect -599 -1908 -433 -1850
rect -341 -1908 -335 -1816
rect -1900 -1914 -335 -1908
rect 335 -1816 439 -1810
rect 335 -1908 341 -1816
rect 433 -1850 439 -1816
rect 593 -1816 697 -1810
rect 593 -1850 599 -1816
rect 433 -1908 599 -1850
rect 691 -1850 697 -1816
rect 1835 -1850 1899 390
rect 691 -1856 1899 -1850
rect 691 -1908 1841 -1856
rect 1893 -1908 1899 -1856
rect 335 -1914 1899 -1908
rect 1999 -1942 2063 2006
rect -2064 -1948 2063 -1942
rect -2064 -2000 -533 -1948
rect -481 -2000 481 -1948
rect 533 -2000 2063 -1948
rect -2064 -2006 2063 -2000
rect 2163 -2034 2227 2190
rect 2487 1976 2551 1982
rect 2487 1924 2493 1976
rect 2545 1924 2551 1976
rect 2487 819 2551 1924
rect 2482 810 2556 819
rect 2482 754 2491 810
rect 2547 754 2556 810
rect 2482 745 2556 754
rect -2228 -2040 2227 -2034
rect -2228 -2092 -1049 -2040
rect -997 -2092 -562 -2040
rect -2228 -2098 -562 -2092
rect -568 -2132 -562 -2098
rect -470 -2092 -26 -2040
rect 26 -2092 470 -2040
rect -470 -2098 470 -2092
rect -470 -2132 -464 -2098
rect -568 -2138 -464 -2132
rect 464 -2132 470 -2098
rect 562 -2092 997 -2040
rect 1049 -2092 2227 -2040
rect 562 -2098 2227 -2092
rect 2327 356 2391 362
rect 2327 304 2333 356
rect 2385 304 2391 356
rect 562 -2132 568 -2098
rect 464 -2138 568 -2132
rect 2327 -2218 2391 304
rect 2487 -360 2551 745
rect 2487 -412 2493 -360
rect 2545 -412 2551 -360
rect 2487 -418 2551 -412
rect -2392 -2282 2391 -2218
rect 2491 -1856 2555 -1850
rect 2491 -1908 2497 -1856
rect 2549 -1908 2555 -1856
rect 2491 -1933 2555 -1908
rect -32 -2310 32 -2282
rect -2096 -2316 2096 -2310
rect -2096 -2368 -2090 -2316
rect -2038 -2368 -1717 -2316
rect -1637 -2368 -1459 -2316
rect -1379 -2368 -1058 -2316
rect -1006 -2368 -427 -2316
rect -347 -2368 -284 -2316
rect -232 -2368 -169 -2316
rect -89 -2368 605 -2316
rect 685 -2368 748 -2316
rect 800 -2368 1006 -2316
rect 1058 -2368 1379 -2316
rect 1459 -2368 1637 -2316
rect 1717 -2368 2038 -2316
rect 2090 -2368 2096 -2316
rect -2096 -2374 2096 -2368
rect -1981 -3632 1981 -3626
rect -1981 -3684 -1975 -3632
rect -1895 -3684 -1574 -3632
rect -1522 -3684 -1201 -3632
rect -1121 -3684 -800 -3632
rect -748 -3684 -685 -3632
rect -605 -3684 89 -3632
rect 169 -3684 232 -3632
rect 284 -3684 347 -3632
rect 427 -3684 1121 -3632
rect 1201 -3684 1522 -3632
rect 1574 -3684 1895 -3632
rect 1975 -3684 1981 -3632
rect -1981 -3690 1981 -3684
rect -32 -3718 32 -3690
rect 2491 -3718 2556 -1933
rect -2556 -3782 2556 -3718
rect -2816 -4016 -2216 -4006
rect -2816 -4326 -2216 -4316
rect 2216 -4016 2816 -4006
rect 2216 -4326 2816 -4316
<< via2 >>
rect -2816 4016 -2216 4316
rect 2216 4016 2816 4316
rect -54 2389 55 2450
rect -966 1955 -910 2011
rect 910 1955 966 2011
rect -1265 514 -1209 570
rect 1199 514 1255 570
rect 2491 754 2547 810
rect -2816 -4316 -2216 -4016
rect 2216 -4316 2816 -4016
<< metal3 >>
rect -2826 4316 -2206 4321
rect -2826 4016 -2816 4316
rect -2216 4016 -2206 4316
rect -2826 4011 -2206 4016
rect 2206 4316 2826 4321
rect 2206 4016 2216 4316
rect 2816 4016 2826 4316
rect 2206 4011 2826 4016
rect -63 2450 63 2459
rect -63 2389 -54 2450
rect 55 2389 63 2450
rect -63 2380 63 2389
rect -2595 2320 63 2380
rect -2595 2153 50 2213
rect -50 2093 50 2153
rect -988 2033 988 2093
rect -988 2011 -888 2033
rect -988 1955 -966 2011
rect -910 1955 -888 2011
rect -988 1933 -888 1955
rect 888 2011 988 2033
rect 888 1955 910 2011
rect 966 1955 988 2011
rect 888 1933 988 1955
rect 2469 812 2569 832
rect 2469 810 2737 812
rect 2469 754 2491 810
rect 2547 754 2737 810
rect 2469 752 2737 754
rect 2469 732 2569 752
rect -1287 570 -1187 592
rect -1287 514 -1265 570
rect -1209 514 -1187 570
rect -1287 492 -1187 514
rect 1177 570 1277 592
rect 1177 514 1199 570
rect 1255 514 1277 570
rect 1177 492 1277 514
rect -1287 432 1277 492
rect -55 372 45 432
rect -2621 312 45 372
rect -2826 -4016 -2206 -4011
rect -2826 -4316 -2816 -4016
rect -2216 -4316 -2206 -4016
rect -2826 -4321 -2206 -4316
rect 2206 -4016 2826 -4011
rect 2206 -4316 2216 -4016
rect 2816 -4316 2826 -4016
rect 2206 -4321 2826 -4316
<< via3 >>
rect -2816 4016 -2216 4316
rect 2216 4016 2816 4316
rect -2816 -4316 -2216 -4016
rect 2216 -4316 2816 -4016
<< metal4 >>
rect -3000 4316 3000 4500
rect -3000 4016 -2816 4316
rect -2216 4016 2216 4316
rect 2816 4016 3000 4316
rect -3000 3700 3000 4016
rect -3000 -4016 3000 -3700
rect -3000 -4316 -2816 -4016
rect -2216 -4316 2216 -4016
rect 2816 -4316 3000 -4016
rect -3000 -4500 3000 -4316
<< labels >>
flabel metal4 -3000 3700 -3000 4500 3 FreeSans 480 0 0 0 vdd
port 2 e
flabel metal3 -2595 2153 -2595 2213 1 FreeSans 280 0 0 0 vinp
port 4 n
flabel metal3 -2621 312 -2621 372 1 FreeSans 280 0 0 0 vinm
port 3 n
flabel metal3 2737 752 2737 812 1 FreeSans 280 0 0 0 vout
port 5 n
flabel metal4 -3000 -4500 -2999 -3700 3 FreeSans 240 0 0 0 vss
port 6 e
flabel metal3 -2595 2320 -2595 2380 1 FreeSans 240 0 0 0 ibias
port 1 n
<< end >>
