magic
tech sky130A
magscale 1 2
timestamp 1624002729
<< error_p >>
rect -1097 566 1097 600
rect -1127 -566 1127 566
rect -1097 -600 1097 -566
<< nwell >>
rect -1097 -600 1097 600
<< mvpmos >>
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
<< mvpdiff >>
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
<< mvpdiffc >>
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
<< poly >>
rect -969 581 -837 597
rect -969 564 -953 581
rect -1003 547 -953 564
rect -853 564 -837 581
rect -711 581 -579 597
rect -711 564 -695 581
rect -853 547 -803 564
rect -1003 500 -803 547
rect -745 547 -695 564
rect -595 564 -579 581
rect -453 581 -321 597
rect -453 564 -437 581
rect -595 547 -545 564
rect -745 500 -545 547
rect -487 547 -437 564
rect -337 564 -321 581
rect -195 581 -63 597
rect -195 564 -179 581
rect -337 547 -287 564
rect -487 500 -287 547
rect -229 547 -179 564
rect -79 564 -63 581
rect 63 581 195 597
rect 63 564 79 581
rect -79 547 -29 564
rect -229 500 -29 547
rect 29 547 79 564
rect 179 564 195 581
rect 321 581 453 597
rect 321 564 337 581
rect 179 547 229 564
rect 29 500 229 547
rect 287 547 337 564
rect 437 564 453 581
rect 579 581 711 597
rect 579 564 595 581
rect 437 547 487 564
rect 287 500 487 547
rect 545 547 595 564
rect 695 564 711 581
rect 837 581 969 597
rect 837 564 853 581
rect 695 547 745 564
rect 545 500 745 547
rect 803 547 853 564
rect 953 564 969 581
rect 953 547 1003 564
rect 803 500 1003 547
rect -1003 -547 -803 -500
rect -1003 -564 -953 -547
rect -969 -581 -953 -564
rect -853 -564 -803 -547
rect -745 -547 -545 -500
rect -745 -564 -695 -547
rect -853 -581 -837 -564
rect -969 -597 -837 -581
rect -711 -581 -695 -564
rect -595 -564 -545 -547
rect -487 -547 -287 -500
rect -487 -564 -437 -547
rect -595 -581 -579 -564
rect -711 -597 -579 -581
rect -453 -581 -437 -564
rect -337 -564 -287 -547
rect -229 -547 -29 -500
rect -229 -564 -179 -547
rect -337 -581 -321 -564
rect -453 -597 -321 -581
rect -195 -581 -179 -564
rect -79 -564 -29 -547
rect 29 -547 229 -500
rect 29 -564 79 -547
rect -79 -581 -63 -564
rect -195 -597 -63 -581
rect 63 -581 79 -564
rect 179 -564 229 -547
rect 287 -547 487 -500
rect 287 -564 337 -547
rect 179 -581 195 -564
rect 63 -597 195 -581
rect 321 -581 337 -564
rect 437 -564 487 -547
rect 545 -547 745 -500
rect 545 -564 595 -547
rect 437 -581 453 -564
rect 321 -597 453 -581
rect 579 -581 595 -564
rect 695 -564 745 -547
rect 803 -547 1003 -500
rect 803 -564 853 -547
rect 695 -581 711 -564
rect 579 -597 711 -581
rect 837 -581 853 -564
rect 953 -564 1003 -547
rect 953 -581 969 -564
rect 837 -597 969 -581
<< polycont >>
rect -953 547 -853 581
rect -695 547 -595 581
rect -437 547 -337 581
rect -179 547 -79 581
rect 79 547 179 581
rect 337 547 437 581
rect 595 547 695 581
rect 853 547 953 581
rect -953 -581 -853 -547
rect -695 -581 -595 -547
rect -437 -581 -337 -547
rect -179 -581 -79 -547
rect 79 -581 179 -547
rect 337 -581 437 -547
rect 595 -581 695 -547
rect 853 -581 953 -547
<< locali >>
rect -969 547 -953 581
rect -853 547 -837 581
rect -711 547 -695 581
rect -595 547 -579 581
rect -453 547 -437 581
rect -337 547 -321 581
rect -195 547 -179 581
rect -79 547 -63 581
rect 63 547 79 581
rect 179 547 195 581
rect 321 547 337 581
rect 437 547 453 581
rect 579 547 595 581
rect 695 547 711 581
rect 837 547 853 581
rect 953 547 969 581
rect -1049 488 -1015 504
rect -1049 -504 -1015 -488
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -504 1049 -488
rect -969 -581 -953 -547
rect -853 -581 -837 -547
rect -711 -581 -695 -547
rect -595 -581 -579 -547
rect -453 -581 -437 -547
rect -337 -581 -321 -547
rect -195 -581 -179 -547
rect -79 -581 -63 -547
rect 63 -581 79 -547
rect 179 -581 195 -547
rect 321 -581 337 -547
rect 437 -581 453 -547
rect 579 -581 595 -547
rect 695 -581 711 -547
rect 837 -581 853 -547
rect 953 -581 969 -547
<< viali >>
rect -937 547 -869 581
rect -679 547 -611 581
rect -421 547 -353 581
rect -163 547 -95 581
rect 95 547 163 581
rect 353 547 421 581
rect 611 547 679 581
rect 869 547 937 581
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect -937 -581 -869 -547
rect -679 -581 -611 -547
rect -421 -581 -353 -547
rect -163 -581 -95 -547
rect 95 -581 163 -547
rect 353 -581 421 -547
rect 611 -581 679 -547
rect 869 -581 937 -547
<< metal1 >>
rect -949 581 -857 587
rect -949 547 -937 581
rect -869 547 -857 581
rect -949 541 -857 547
rect -691 581 -599 587
rect -691 547 -679 581
rect -611 547 -599 581
rect -691 541 -599 547
rect -433 581 -341 587
rect -433 547 -421 581
rect -353 547 -341 581
rect -433 541 -341 547
rect -175 581 -83 587
rect -175 547 -163 581
rect -95 547 -83 581
rect -175 541 -83 547
rect 83 581 175 587
rect 83 547 95 581
rect 163 547 175 581
rect 83 541 175 547
rect 341 581 433 587
rect 341 547 353 581
rect 421 547 433 581
rect 341 541 433 547
rect 599 581 691 587
rect 599 547 611 581
rect 679 547 691 581
rect 599 541 691 547
rect 857 581 949 587
rect 857 547 869 581
rect 937 547 949 581
rect 857 541 949 547
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect -949 -547 -857 -541
rect -949 -581 -937 -547
rect -869 -581 -857 -547
rect -949 -587 -857 -581
rect -691 -547 -599 -541
rect -691 -581 -679 -547
rect -611 -581 -599 -547
rect -691 -587 -599 -581
rect -433 -547 -341 -541
rect -433 -581 -421 -547
rect -353 -581 -341 -547
rect -433 -587 -341 -581
rect -175 -547 -83 -541
rect -175 -581 -163 -547
rect -95 -581 -83 -547
rect -175 -587 -83 -581
rect 83 -547 175 -541
rect 83 -581 95 -547
rect 163 -581 175 -547
rect 83 -587 175 -581
rect 341 -547 433 -541
rect 341 -581 353 -547
rect 421 -581 433 -547
rect 341 -587 433 -581
rect 599 -547 691 -541
rect 599 -581 611 -547
rect 679 -581 691 -547
rect 599 -587 691 -581
rect 857 -547 949 -541
rect 857 -581 869 -547
rect 937 -581 949 -547
rect 857 -587 949 -581
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string parameters w 5 l 1 m 1 nf 8 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
