magic
tech sky130A
magscale 1 2
timestamp 1624002729
<< poly >>
rect -200 687 200 703
rect -200 653 -184 687
rect 184 653 200 687
rect -200 630 200 653
rect -200 -653 200 -630
rect -200 -687 -184 -653
rect 184 -687 200 -653
rect -200 -703 200 -687
<< polycont >>
rect -184 653 184 687
rect -184 -687 184 -653
<< npolyres >>
rect -200 -630 200 630
<< locali >>
rect -200 653 -184 687
rect 184 653 200 687
rect -200 -687 -184 -653
rect 184 -687 200 -653
<< viali >>
rect -184 653 184 687
rect -184 647 184 653
rect -184 -653 184 -647
rect -184 -687 184 -653
<< metal1 >>
rect -196 687 196 693
rect -196 647 -184 687
rect 184 647 196 687
rect -196 641 196 647
rect -196 -647 196 -641
rect -196 -687 -184 -647
rect 184 -687 196 -647
rect -196 -693 196 -687
<< properties >>
string gencell sky130_fd_pr__res_generic_po
string parameters w 2 l 6.3 m 1 nx 1 wmin 0.330 lmin 1.650 rho 48.2 val 151.83 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
