magic
tech sky130A
magscale 1 2
timestamp 1624002729
<< dnwell >>
rect -2300 -3300 2300 -740
<< nwell >>
rect -2000 400 2000 2400
rect -2400 -1000 2400 -640
rect -2400 -3000 -2000 -1000
rect 2000 -3000 2400 -1000
rect -2400 -3400 2400 -3000
<< pwell >>
rect -2400 2400 2400 2800
rect -2400 400 -2000 2400
rect 2000 400 2400 2400
rect -2400 40 2400 400
rect -2000 -3000 2000 -1000
<< mvnmos >>
rect -1551 -2500 -1451 -1500
rect -1393 -2500 -1293 -1500
rect -1235 -2500 -1135 -1500
rect -1077 -2500 -977 -1500
rect -919 -2500 -819 -1500
rect -761 -2500 -661 -1500
rect -603 -2500 -503 -1500
rect -445 -2500 -345 -1500
rect -287 -2500 -187 -1500
rect -129 -2500 -29 -1500
rect 29 -2500 129 -1500
rect 187 -2500 287 -1500
rect 345 -2500 445 -1500
rect 503 -2500 603 -1500
rect 661 -2500 761 -1500
rect 819 -2500 919 -1500
rect 977 -2500 1077 -1500
rect 1135 -2500 1235 -1500
rect 1293 -2500 1393 -1500
rect 1451 -2500 1551 -1500
<< mvpmos >>
rect -1551 900 -1451 1900
rect -1393 900 -1293 1900
rect -1235 900 -1135 1900
rect -1077 900 -977 1900
rect -919 900 -819 1900
rect -761 900 -661 1900
rect -603 900 -503 1900
rect -445 900 -345 1900
rect -287 900 -187 1900
rect -129 900 -29 1900
rect 29 900 129 1900
rect 187 900 287 1900
rect 345 900 445 1900
rect 503 900 603 1900
rect 661 900 761 1900
rect 819 900 919 1900
rect 977 900 1077 1900
rect 1135 900 1235 1900
rect 1293 900 1393 1900
rect 1451 900 1551 1900
<< mvndiff >>
rect -1609 -1512 -1551 -1500
rect -1609 -2488 -1597 -1512
rect -1563 -2488 -1551 -1512
rect -1609 -2500 -1551 -2488
rect -1451 -1512 -1393 -1500
rect -1451 -2488 -1439 -1512
rect -1405 -2488 -1393 -1512
rect -1451 -2500 -1393 -2488
rect -1293 -1512 -1235 -1500
rect -1293 -2488 -1281 -1512
rect -1247 -2488 -1235 -1512
rect -1293 -2500 -1235 -2488
rect -1135 -1512 -1077 -1500
rect -1135 -2488 -1123 -1512
rect -1089 -2488 -1077 -1512
rect -1135 -2500 -1077 -2488
rect -977 -1512 -919 -1500
rect -977 -2488 -965 -1512
rect -931 -2488 -919 -1512
rect -977 -2500 -919 -2488
rect -819 -1512 -761 -1500
rect -819 -2488 -807 -1512
rect -773 -2488 -761 -1512
rect -819 -2500 -761 -2488
rect -661 -1512 -603 -1500
rect -661 -2488 -649 -1512
rect -615 -2488 -603 -1512
rect -661 -2500 -603 -2488
rect -503 -1512 -445 -1500
rect -503 -2488 -491 -1512
rect -457 -2488 -445 -1512
rect -503 -2500 -445 -2488
rect -345 -1512 -287 -1500
rect -345 -2488 -333 -1512
rect -299 -2488 -287 -1512
rect -345 -2500 -287 -2488
rect -187 -1512 -129 -1500
rect -187 -2488 -175 -1512
rect -141 -2488 -129 -1512
rect -187 -2500 -129 -2488
rect -29 -1512 29 -1500
rect -29 -2488 -17 -1512
rect 17 -2488 29 -1512
rect -29 -2500 29 -2488
rect 129 -1512 187 -1500
rect 129 -2488 141 -1512
rect 175 -2488 187 -1512
rect 129 -2500 187 -2488
rect 287 -1512 345 -1500
rect 287 -2488 299 -1512
rect 333 -2488 345 -1512
rect 287 -2500 345 -2488
rect 445 -1512 503 -1500
rect 445 -2488 457 -1512
rect 491 -2488 503 -1512
rect 445 -2500 503 -2488
rect 603 -1512 661 -1500
rect 603 -2488 615 -1512
rect 649 -2488 661 -1512
rect 603 -2500 661 -2488
rect 761 -1512 819 -1500
rect 761 -2488 773 -1512
rect 807 -2488 819 -1512
rect 761 -2500 819 -2488
rect 919 -1512 977 -1500
rect 919 -2488 931 -1512
rect 965 -2488 977 -1512
rect 919 -2500 977 -2488
rect 1077 -1512 1135 -1500
rect 1077 -2488 1089 -1512
rect 1123 -2488 1135 -1512
rect 1077 -2500 1135 -2488
rect 1235 -1512 1293 -1500
rect 1235 -2488 1247 -1512
rect 1281 -2488 1293 -1512
rect 1235 -2500 1293 -2488
rect 1393 -1512 1451 -1500
rect 1393 -2488 1405 -1512
rect 1439 -2488 1451 -1512
rect 1393 -2500 1451 -2488
rect 1551 -1512 1609 -1500
rect 1551 -2488 1563 -1512
rect 1597 -2488 1609 -1512
rect 1551 -2500 1609 -2488
<< mvpdiff >>
rect -1609 1888 -1551 1900
rect -1609 912 -1597 1888
rect -1563 912 -1551 1888
rect -1609 900 -1551 912
rect -1451 1888 -1393 1900
rect -1451 912 -1439 1888
rect -1405 912 -1393 1888
rect -1451 900 -1393 912
rect -1293 1888 -1235 1900
rect -1293 912 -1281 1888
rect -1247 912 -1235 1888
rect -1293 900 -1235 912
rect -1135 1888 -1077 1900
rect -1135 912 -1123 1888
rect -1089 912 -1077 1888
rect -1135 900 -1077 912
rect -977 1888 -919 1900
rect -977 912 -965 1888
rect -931 912 -919 1888
rect -977 900 -919 912
rect -819 1888 -761 1900
rect -819 912 -807 1888
rect -773 912 -761 1888
rect -819 900 -761 912
rect -661 1888 -603 1900
rect -661 912 -649 1888
rect -615 912 -603 1888
rect -661 900 -603 912
rect -503 1888 -445 1900
rect -503 912 -491 1888
rect -457 912 -445 1888
rect -503 900 -445 912
rect -345 1888 -287 1900
rect -345 912 -333 1888
rect -299 912 -287 1888
rect -345 900 -287 912
rect -187 1888 -129 1900
rect -187 912 -175 1888
rect -141 912 -129 1888
rect -187 900 -129 912
rect -29 1888 29 1900
rect -29 912 -17 1888
rect 17 912 29 1888
rect -29 900 29 912
rect 129 1888 187 1900
rect 129 912 141 1888
rect 175 912 187 1888
rect 129 900 187 912
rect 287 1888 345 1900
rect 287 912 299 1888
rect 333 912 345 1888
rect 287 900 345 912
rect 445 1888 503 1900
rect 445 912 457 1888
rect 491 912 503 1888
rect 445 900 503 912
rect 603 1888 661 1900
rect 603 912 615 1888
rect 649 912 661 1888
rect 603 900 661 912
rect 761 1888 819 1900
rect 761 912 773 1888
rect 807 912 819 1888
rect 761 900 819 912
rect 919 1888 977 1900
rect 919 912 931 1888
rect 965 912 977 1888
rect 919 900 977 912
rect 1077 1888 1135 1900
rect 1077 912 1089 1888
rect 1123 912 1135 1888
rect 1077 900 1135 912
rect 1235 1888 1293 1900
rect 1235 912 1247 1888
rect 1281 912 1293 1888
rect 1235 900 1293 912
rect 1393 1888 1451 1900
rect 1393 912 1405 1888
rect 1439 912 1451 1888
rect 1393 900 1451 912
rect 1551 1888 1609 1900
rect 1551 912 1563 1888
rect 1597 912 1609 1888
rect 1551 900 1609 912
<< mvndiffc >>
rect -1597 -2488 -1563 -1512
rect -1439 -2488 -1405 -1512
rect -1281 -2488 -1247 -1512
rect -1123 -2488 -1089 -1512
rect -965 -2488 -931 -1512
rect -807 -2488 -773 -1512
rect -649 -2488 -615 -1512
rect -491 -2488 -457 -1512
rect -333 -2488 -299 -1512
rect -175 -2488 -141 -1512
rect -17 -2488 17 -1512
rect 141 -2488 175 -1512
rect 299 -2488 333 -1512
rect 457 -2488 491 -1512
rect 615 -2488 649 -1512
rect 773 -2488 807 -1512
rect 931 -2488 965 -1512
rect 1089 -2488 1123 -1512
rect 1247 -2488 1281 -1512
rect 1405 -2488 1439 -1512
rect 1563 -2488 1597 -1512
<< mvpdiffc >>
rect -1597 912 -1563 1888
rect -1439 912 -1405 1888
rect -1281 912 -1247 1888
rect -1123 912 -1089 1888
rect -965 912 -931 1888
rect -807 912 -773 1888
rect -649 912 -615 1888
rect -491 912 -457 1888
rect -333 912 -299 1888
rect -175 912 -141 1888
rect -17 912 17 1888
rect 141 912 175 1888
rect 299 912 333 1888
rect 457 912 491 1888
rect 615 912 649 1888
rect 773 912 807 1888
rect 931 912 965 1888
rect 1089 912 1123 1888
rect 1247 912 1281 1888
rect 1405 912 1439 1888
rect 1563 912 1597 1888
<< mvpsubdiff >>
rect -2334 2722 2334 2734
rect -2334 2562 -2100 2722
rect 2100 2562 2334 2722
rect -2334 2550 2334 2562
rect -2334 2500 -2150 2550
rect -2334 340 -2322 2500
rect -2162 340 -2150 2500
rect 2150 2500 2334 2550
rect -2334 290 -2150 340
rect 2150 340 2162 2500
rect 2322 340 2334 2500
rect 2150 290 2334 340
rect -2334 278 2334 290
rect -2334 118 -2100 278
rect 2100 118 2334 278
rect -2334 106 2334 118
rect -1934 -1078 1934 -1066
rect -1934 -1238 -1700 -1078
rect 1700 -1238 1934 -1078
rect -1934 -1250 1934 -1238
rect -1934 -1300 -1750 -1250
rect -1934 -2700 -1922 -1300
rect -1762 -2700 -1750 -1300
rect 1750 -1300 1934 -1250
rect -1934 -2750 -1750 -2700
rect 1750 -2700 1762 -1300
rect 1922 -2700 1934 -1300
rect 1750 -2750 1934 -2700
rect -1934 -2762 1934 -2750
rect -1934 -2922 -1700 -2762
rect 1700 -2922 1934 -2762
rect -1934 -2934 1934 -2922
<< mvnsubdiff >>
rect -1934 2322 1934 2334
rect -1934 2162 -1700 2322
rect 1700 2162 1934 2322
rect -1934 2150 1934 2162
rect -1934 2100 -1750 2150
rect -1934 700 -1922 2100
rect -1762 700 -1750 2100
rect 1750 2100 1934 2150
rect -1934 650 -1750 700
rect 1750 700 1762 2100
rect 1922 700 1934 2100
rect 1750 650 1934 700
rect -1934 638 1934 650
rect -1934 478 -1700 638
rect 1700 478 1934 638
rect -1934 466 1934 478
rect -2334 -718 2334 -706
rect -2334 -878 -2100 -718
rect 2100 -878 2334 -718
rect -2334 -890 2334 -878
rect -2334 -940 -2150 -890
rect -2334 -3100 -2322 -940
rect -2162 -3100 -2150 -940
rect 2150 -940 2334 -890
rect -2334 -3150 -2150 -3100
rect 2150 -3100 2162 -940
rect 2322 -3100 2334 -940
rect 2150 -3150 2334 -3100
rect -2334 -3162 2334 -3150
rect -2334 -3322 -2100 -3162
rect 2100 -3322 2334 -3162
rect -2334 -3334 2334 -3322
<< mvpsubdiffcont >>
rect -2100 2562 2100 2722
rect -2322 340 -2162 2500
rect 2162 340 2322 2500
rect -2100 118 2100 278
rect -1700 -1238 1700 -1078
rect -1922 -2700 -1762 -1300
rect 1762 -2700 1922 -1300
rect -1700 -2922 1700 -2762
<< mvnsubdiffcont >>
rect -1700 2162 1700 2322
rect -1922 700 -1762 2100
rect 1762 700 1922 2100
rect -1700 478 1700 638
rect -2100 -878 2100 -718
rect -2322 -3100 -2162 -940
rect 2162 -3100 2322 -940
rect -2100 -3322 2100 -3162
<< poly >>
rect -1537 1981 -1465 1997
rect -1537 1964 -1521 1981
rect -1551 1947 -1521 1964
rect -1481 1964 -1465 1981
rect -1379 1981 -1307 1997
rect -1379 1964 -1363 1981
rect -1481 1947 -1451 1964
rect -1551 1900 -1451 1947
rect -1393 1947 -1363 1964
rect -1323 1964 -1307 1981
rect -1221 1981 -1149 1997
rect -1221 1964 -1205 1981
rect -1323 1947 -1293 1964
rect -1393 1900 -1293 1947
rect -1235 1947 -1205 1964
rect -1165 1964 -1149 1981
rect -1063 1981 -991 1997
rect -1063 1964 -1047 1981
rect -1165 1947 -1135 1964
rect -1235 1900 -1135 1947
rect -1077 1947 -1047 1964
rect -1007 1964 -991 1981
rect -905 1981 -833 1997
rect -905 1964 -889 1981
rect -1007 1947 -977 1964
rect -1077 1900 -977 1947
rect -919 1947 -889 1964
rect -849 1964 -833 1981
rect -747 1981 -675 1997
rect -747 1964 -731 1981
rect -849 1947 -819 1964
rect -919 1900 -819 1947
rect -761 1947 -731 1964
rect -691 1964 -675 1981
rect -589 1981 -517 1997
rect -589 1964 -573 1981
rect -691 1947 -661 1964
rect -761 1900 -661 1947
rect -603 1947 -573 1964
rect -533 1964 -517 1981
rect -431 1981 -359 1997
rect -431 1964 -415 1981
rect -533 1947 -503 1964
rect -603 1900 -503 1947
rect -445 1947 -415 1964
rect -375 1964 -359 1981
rect -273 1981 -201 1997
rect -273 1964 -257 1981
rect -375 1947 -345 1964
rect -445 1900 -345 1947
rect -287 1947 -257 1964
rect -217 1964 -201 1981
rect -115 1981 -43 1997
rect -115 1964 -99 1981
rect -217 1947 -187 1964
rect -287 1900 -187 1947
rect -129 1947 -99 1964
rect -59 1964 -43 1981
rect 43 1981 115 1997
rect 43 1964 59 1981
rect -59 1947 -29 1964
rect -129 1900 -29 1947
rect 29 1947 59 1964
rect 99 1964 115 1981
rect 201 1981 273 1997
rect 201 1964 217 1981
rect 99 1947 129 1964
rect 29 1900 129 1947
rect 187 1947 217 1964
rect 257 1964 273 1981
rect 359 1981 431 1997
rect 359 1964 375 1981
rect 257 1947 287 1964
rect 187 1900 287 1947
rect 345 1947 375 1964
rect 415 1964 431 1981
rect 517 1981 589 1997
rect 517 1964 533 1981
rect 415 1947 445 1964
rect 345 1900 445 1947
rect 503 1947 533 1964
rect 573 1964 589 1981
rect 675 1981 747 1997
rect 675 1964 691 1981
rect 573 1947 603 1964
rect 503 1900 603 1947
rect 661 1947 691 1964
rect 731 1964 747 1981
rect 833 1981 905 1997
rect 833 1964 849 1981
rect 731 1947 761 1964
rect 661 1900 761 1947
rect 819 1947 849 1964
rect 889 1964 905 1981
rect 991 1981 1063 1997
rect 991 1964 1007 1981
rect 889 1947 919 1964
rect 819 1900 919 1947
rect 977 1947 1007 1964
rect 1047 1964 1063 1981
rect 1149 1981 1221 1997
rect 1149 1964 1165 1981
rect 1047 1947 1077 1964
rect 977 1900 1077 1947
rect 1135 1947 1165 1964
rect 1205 1964 1221 1981
rect 1307 1981 1379 1997
rect 1307 1964 1323 1981
rect 1205 1947 1235 1964
rect 1135 1900 1235 1947
rect 1293 1947 1323 1964
rect 1363 1964 1379 1981
rect 1465 1981 1537 1997
rect 1465 1964 1481 1981
rect 1363 1947 1393 1964
rect 1293 1900 1393 1947
rect 1451 1947 1481 1964
rect 1521 1964 1537 1981
rect 1521 1947 1551 1964
rect 1451 1900 1551 1947
rect -1551 853 -1451 900
rect -1551 836 -1521 853
rect -1537 819 -1521 836
rect -1481 836 -1451 853
rect -1393 853 -1293 900
rect -1393 836 -1363 853
rect -1481 819 -1465 836
rect -1537 803 -1465 819
rect -1379 819 -1363 836
rect -1323 836 -1293 853
rect -1235 853 -1135 900
rect -1235 836 -1205 853
rect -1323 819 -1307 836
rect -1379 803 -1307 819
rect -1221 819 -1205 836
rect -1165 836 -1135 853
rect -1077 853 -977 900
rect -1077 836 -1047 853
rect -1165 819 -1149 836
rect -1221 803 -1149 819
rect -1063 819 -1047 836
rect -1007 836 -977 853
rect -919 853 -819 900
rect -919 836 -889 853
rect -1007 819 -991 836
rect -1063 803 -991 819
rect -905 819 -889 836
rect -849 836 -819 853
rect -761 853 -661 900
rect -761 836 -731 853
rect -849 819 -833 836
rect -905 803 -833 819
rect -747 819 -731 836
rect -691 836 -661 853
rect -603 853 -503 900
rect -603 836 -573 853
rect -691 819 -675 836
rect -747 803 -675 819
rect -589 819 -573 836
rect -533 836 -503 853
rect -445 853 -345 900
rect -445 836 -415 853
rect -533 819 -517 836
rect -589 803 -517 819
rect -431 819 -415 836
rect -375 836 -345 853
rect -287 853 -187 900
rect -287 836 -257 853
rect -375 819 -359 836
rect -431 803 -359 819
rect -273 819 -257 836
rect -217 836 -187 853
rect -129 853 -29 900
rect -129 836 -99 853
rect -217 819 -201 836
rect -273 803 -201 819
rect -115 819 -99 836
rect -59 836 -29 853
rect 29 853 129 900
rect 29 836 59 853
rect -59 819 -43 836
rect -115 803 -43 819
rect 43 819 59 836
rect 99 836 129 853
rect 187 853 287 900
rect 187 836 217 853
rect 99 819 115 836
rect 43 803 115 819
rect 201 819 217 836
rect 257 836 287 853
rect 345 853 445 900
rect 345 836 375 853
rect 257 819 273 836
rect 201 803 273 819
rect 359 819 375 836
rect 415 836 445 853
rect 503 853 603 900
rect 503 836 533 853
rect 415 819 431 836
rect 359 803 431 819
rect 517 819 533 836
rect 573 836 603 853
rect 661 853 761 900
rect 661 836 691 853
rect 573 819 589 836
rect 517 803 589 819
rect 675 819 691 836
rect 731 836 761 853
rect 819 853 919 900
rect 819 836 849 853
rect 731 819 747 836
rect 675 803 747 819
rect 833 819 849 836
rect 889 836 919 853
rect 977 853 1077 900
rect 977 836 1007 853
rect 889 819 905 836
rect 833 803 905 819
rect 991 819 1007 836
rect 1047 836 1077 853
rect 1135 853 1235 900
rect 1135 836 1165 853
rect 1047 819 1063 836
rect 991 803 1063 819
rect 1149 819 1165 836
rect 1205 836 1235 853
rect 1293 853 1393 900
rect 1293 836 1323 853
rect 1205 819 1221 836
rect 1149 803 1221 819
rect 1307 819 1323 836
rect 1363 836 1393 853
rect 1451 853 1551 900
rect 1451 836 1481 853
rect 1363 819 1379 836
rect 1307 803 1379 819
rect 1465 819 1481 836
rect 1521 836 1551 853
rect 1521 819 1537 836
rect 1465 803 1537 819
rect -1537 -1428 -1465 -1412
rect -1537 -1445 -1521 -1428
rect -1551 -1462 -1521 -1445
rect -1481 -1445 -1465 -1428
rect -1379 -1428 -1307 -1412
rect -1379 -1445 -1363 -1428
rect -1481 -1462 -1451 -1445
rect -1551 -1500 -1451 -1462
rect -1393 -1462 -1363 -1445
rect -1323 -1445 -1307 -1428
rect -1221 -1428 -1149 -1412
rect -1221 -1445 -1205 -1428
rect -1323 -1462 -1293 -1445
rect -1393 -1500 -1293 -1462
rect -1235 -1462 -1205 -1445
rect -1165 -1445 -1149 -1428
rect -1063 -1428 -991 -1412
rect -1063 -1445 -1047 -1428
rect -1165 -1462 -1135 -1445
rect -1235 -1500 -1135 -1462
rect -1077 -1462 -1047 -1445
rect -1007 -1445 -991 -1428
rect -905 -1428 -833 -1412
rect -905 -1445 -889 -1428
rect -1007 -1462 -977 -1445
rect -1077 -1500 -977 -1462
rect -919 -1462 -889 -1445
rect -849 -1445 -833 -1428
rect -747 -1428 -675 -1412
rect -747 -1445 -731 -1428
rect -849 -1462 -819 -1445
rect -919 -1500 -819 -1462
rect -761 -1462 -731 -1445
rect -691 -1445 -675 -1428
rect -589 -1428 -517 -1412
rect -589 -1445 -573 -1428
rect -691 -1462 -661 -1445
rect -761 -1500 -661 -1462
rect -603 -1462 -573 -1445
rect -533 -1445 -517 -1428
rect -431 -1428 -359 -1412
rect -431 -1445 -415 -1428
rect -533 -1462 -503 -1445
rect -603 -1500 -503 -1462
rect -445 -1462 -415 -1445
rect -375 -1445 -359 -1428
rect -273 -1428 -201 -1412
rect -273 -1445 -257 -1428
rect -375 -1462 -345 -1445
rect -445 -1500 -345 -1462
rect -287 -1462 -257 -1445
rect -217 -1445 -201 -1428
rect -115 -1428 -43 -1412
rect -115 -1445 -99 -1428
rect -217 -1462 -187 -1445
rect -287 -1500 -187 -1462
rect -129 -1462 -99 -1445
rect -59 -1445 -43 -1428
rect 43 -1428 115 -1412
rect 43 -1445 59 -1428
rect -59 -1462 -29 -1445
rect -129 -1500 -29 -1462
rect 29 -1462 59 -1445
rect 99 -1445 115 -1428
rect 201 -1428 273 -1412
rect 201 -1445 217 -1428
rect 99 -1462 129 -1445
rect 29 -1500 129 -1462
rect 187 -1462 217 -1445
rect 257 -1445 273 -1428
rect 359 -1428 431 -1412
rect 359 -1445 375 -1428
rect 257 -1462 287 -1445
rect 187 -1500 287 -1462
rect 345 -1462 375 -1445
rect 415 -1445 431 -1428
rect 517 -1428 589 -1412
rect 517 -1445 533 -1428
rect 415 -1462 445 -1445
rect 345 -1500 445 -1462
rect 503 -1462 533 -1445
rect 573 -1445 589 -1428
rect 675 -1428 747 -1412
rect 675 -1445 691 -1428
rect 573 -1462 603 -1445
rect 503 -1500 603 -1462
rect 661 -1462 691 -1445
rect 731 -1445 747 -1428
rect 833 -1428 905 -1412
rect 833 -1445 849 -1428
rect 731 -1462 761 -1445
rect 661 -1500 761 -1462
rect 819 -1462 849 -1445
rect 889 -1445 905 -1428
rect 991 -1428 1063 -1412
rect 991 -1445 1007 -1428
rect 889 -1462 919 -1445
rect 819 -1500 919 -1462
rect 977 -1462 1007 -1445
rect 1047 -1445 1063 -1428
rect 1149 -1428 1221 -1412
rect 1149 -1445 1165 -1428
rect 1047 -1462 1077 -1445
rect 977 -1500 1077 -1462
rect 1135 -1462 1165 -1445
rect 1205 -1445 1221 -1428
rect 1307 -1428 1379 -1412
rect 1307 -1445 1323 -1428
rect 1205 -1462 1235 -1445
rect 1135 -1500 1235 -1462
rect 1293 -1462 1323 -1445
rect 1363 -1445 1379 -1428
rect 1465 -1428 1537 -1412
rect 1465 -1445 1481 -1428
rect 1363 -1462 1393 -1445
rect 1293 -1500 1393 -1462
rect 1451 -1462 1481 -1445
rect 1521 -1445 1537 -1428
rect 1521 -1462 1551 -1445
rect 1451 -1500 1551 -1462
rect -1551 -2538 -1451 -2500
rect -1551 -2555 -1521 -2538
rect -1537 -2572 -1521 -2555
rect -1481 -2555 -1451 -2538
rect -1393 -2538 -1293 -2500
rect -1393 -2555 -1363 -2538
rect -1481 -2572 -1465 -2555
rect -1537 -2588 -1465 -2572
rect -1379 -2572 -1363 -2555
rect -1323 -2555 -1293 -2538
rect -1235 -2538 -1135 -2500
rect -1235 -2555 -1205 -2538
rect -1323 -2572 -1307 -2555
rect -1379 -2588 -1307 -2572
rect -1221 -2572 -1205 -2555
rect -1165 -2555 -1135 -2538
rect -1077 -2538 -977 -2500
rect -1077 -2555 -1047 -2538
rect -1165 -2572 -1149 -2555
rect -1221 -2588 -1149 -2572
rect -1063 -2572 -1047 -2555
rect -1007 -2555 -977 -2538
rect -919 -2538 -819 -2500
rect -919 -2555 -889 -2538
rect -1007 -2572 -991 -2555
rect -1063 -2588 -991 -2572
rect -905 -2572 -889 -2555
rect -849 -2555 -819 -2538
rect -761 -2538 -661 -2500
rect -761 -2555 -731 -2538
rect -849 -2572 -833 -2555
rect -905 -2588 -833 -2572
rect -747 -2572 -731 -2555
rect -691 -2555 -661 -2538
rect -603 -2538 -503 -2500
rect -603 -2555 -573 -2538
rect -691 -2572 -675 -2555
rect -747 -2588 -675 -2572
rect -589 -2572 -573 -2555
rect -533 -2555 -503 -2538
rect -445 -2538 -345 -2500
rect -445 -2555 -415 -2538
rect -533 -2572 -517 -2555
rect -589 -2588 -517 -2572
rect -431 -2572 -415 -2555
rect -375 -2555 -345 -2538
rect -287 -2538 -187 -2500
rect -287 -2555 -257 -2538
rect -375 -2572 -359 -2555
rect -431 -2588 -359 -2572
rect -273 -2572 -257 -2555
rect -217 -2555 -187 -2538
rect -129 -2538 -29 -2500
rect -129 -2555 -99 -2538
rect -217 -2572 -201 -2555
rect -273 -2588 -201 -2572
rect -115 -2572 -99 -2555
rect -59 -2555 -29 -2538
rect 29 -2538 129 -2500
rect 29 -2555 59 -2538
rect -59 -2572 -43 -2555
rect -115 -2588 -43 -2572
rect 43 -2572 59 -2555
rect 99 -2555 129 -2538
rect 187 -2538 287 -2500
rect 187 -2555 217 -2538
rect 99 -2572 115 -2555
rect 43 -2588 115 -2572
rect 201 -2572 217 -2555
rect 257 -2555 287 -2538
rect 345 -2538 445 -2500
rect 345 -2555 375 -2538
rect 257 -2572 273 -2555
rect 201 -2588 273 -2572
rect 359 -2572 375 -2555
rect 415 -2555 445 -2538
rect 503 -2538 603 -2500
rect 503 -2555 533 -2538
rect 415 -2572 431 -2555
rect 359 -2588 431 -2572
rect 517 -2572 533 -2555
rect 573 -2555 603 -2538
rect 661 -2538 761 -2500
rect 661 -2555 691 -2538
rect 573 -2572 589 -2555
rect 517 -2588 589 -2572
rect 675 -2572 691 -2555
rect 731 -2555 761 -2538
rect 819 -2538 919 -2500
rect 819 -2555 849 -2538
rect 731 -2572 747 -2555
rect 675 -2588 747 -2572
rect 833 -2572 849 -2555
rect 889 -2555 919 -2538
rect 977 -2538 1077 -2500
rect 977 -2555 1007 -2538
rect 889 -2572 905 -2555
rect 833 -2588 905 -2572
rect 991 -2572 1007 -2555
rect 1047 -2555 1077 -2538
rect 1135 -2538 1235 -2500
rect 1135 -2555 1165 -2538
rect 1047 -2572 1063 -2555
rect 991 -2588 1063 -2572
rect 1149 -2572 1165 -2555
rect 1205 -2555 1235 -2538
rect 1293 -2538 1393 -2500
rect 1293 -2555 1323 -2538
rect 1205 -2572 1221 -2555
rect 1149 -2588 1221 -2572
rect 1307 -2572 1323 -2555
rect 1363 -2555 1393 -2538
rect 1451 -2538 1551 -2500
rect 1451 -2555 1481 -2538
rect 1363 -2572 1379 -2555
rect 1307 -2588 1379 -2572
rect 1465 -2572 1481 -2555
rect 1521 -2555 1551 -2538
rect 1521 -2572 1537 -2555
rect 1465 -2588 1537 -2572
<< polycont >>
rect -1521 1947 -1481 1981
rect -1363 1947 -1323 1981
rect -1205 1947 -1165 1981
rect -1047 1947 -1007 1981
rect -889 1947 -849 1981
rect -731 1947 -691 1981
rect -573 1947 -533 1981
rect -415 1947 -375 1981
rect -257 1947 -217 1981
rect -99 1947 -59 1981
rect 59 1947 99 1981
rect 217 1947 257 1981
rect 375 1947 415 1981
rect 533 1947 573 1981
rect 691 1947 731 1981
rect 849 1947 889 1981
rect 1007 1947 1047 1981
rect 1165 1947 1205 1981
rect 1323 1947 1363 1981
rect 1481 1947 1521 1981
rect -1521 819 -1481 853
rect -1363 819 -1323 853
rect -1205 819 -1165 853
rect -1047 819 -1007 853
rect -889 819 -849 853
rect -731 819 -691 853
rect -573 819 -533 853
rect -415 819 -375 853
rect -257 819 -217 853
rect -99 819 -59 853
rect 59 819 99 853
rect 217 819 257 853
rect 375 819 415 853
rect 533 819 573 853
rect 691 819 731 853
rect 849 819 889 853
rect 1007 819 1047 853
rect 1165 819 1205 853
rect 1323 819 1363 853
rect 1481 819 1521 853
rect -1521 -1462 -1481 -1428
rect -1363 -1462 -1323 -1428
rect -1205 -1462 -1165 -1428
rect -1047 -1462 -1007 -1428
rect -889 -1462 -849 -1428
rect -731 -1462 -691 -1428
rect -573 -1462 -533 -1428
rect -415 -1462 -375 -1428
rect -257 -1462 -217 -1428
rect -99 -1462 -59 -1428
rect 59 -1462 99 -1428
rect 217 -1462 257 -1428
rect 375 -1462 415 -1428
rect 533 -1462 573 -1428
rect 691 -1462 731 -1428
rect 849 -1462 889 -1428
rect 1007 -1462 1047 -1428
rect 1165 -1462 1205 -1428
rect 1323 -1462 1363 -1428
rect 1481 -1462 1521 -1428
rect -1521 -2572 -1481 -2538
rect -1363 -2572 -1323 -2538
rect -1205 -2572 -1165 -2538
rect -1047 -2572 -1007 -2538
rect -889 -2572 -849 -2538
rect -731 -2572 -691 -2538
rect -573 -2572 -533 -2538
rect -415 -2572 -375 -2538
rect -257 -2572 -217 -2538
rect -99 -2572 -59 -2538
rect 59 -2572 99 -2538
rect 217 -2572 257 -2538
rect 375 -2572 415 -2538
rect 533 -2572 573 -2538
rect 691 -2572 731 -2538
rect 849 -2572 889 -2538
rect 1007 -2572 1047 -2538
rect 1165 -2572 1205 -2538
rect 1323 -2572 1363 -2538
rect 1481 -2572 1521 -2538
<< locali >>
rect -2322 2500 -2162 2722
rect 2162 2500 2322 2722
rect -1922 2100 -1762 2322
rect 1762 2100 1922 2322
rect -1597 1888 -1563 1904
rect -1597 896 -1563 912
rect -1439 1888 -1405 1904
rect -1439 896 -1405 912
rect -1281 1888 -1247 1904
rect -1281 896 -1247 912
rect -1123 1888 -1089 1904
rect -1123 896 -1089 912
rect -965 1888 -931 1904
rect -965 896 -931 912
rect -807 1888 -773 1904
rect -807 896 -773 912
rect -649 1888 -615 1904
rect -649 896 -615 912
rect -491 1888 -457 1904
rect -491 896 -457 912
rect -333 1888 -299 1904
rect -333 896 -299 912
rect -175 1888 -141 1904
rect -175 896 -141 912
rect -17 1888 17 1904
rect -17 896 17 912
rect 141 1888 175 1904
rect 141 896 175 912
rect 299 1888 333 1904
rect 299 896 333 912
rect 457 1888 491 1904
rect 457 896 491 912
rect 615 1888 649 1904
rect 615 896 649 912
rect 773 1888 807 1904
rect 773 896 807 912
rect 931 1888 965 1904
rect 931 896 965 912
rect 1089 1888 1123 1904
rect 1089 896 1123 912
rect 1247 1888 1281 1904
rect 1247 896 1281 912
rect 1405 1888 1439 1904
rect 1405 896 1439 912
rect 1563 1888 1597 1904
rect 1563 896 1597 912
rect -1537 819 -1521 853
rect -1481 819 -1465 853
rect -1379 819 -1363 853
rect -1323 819 -1307 853
rect -1221 819 -1205 853
rect -1165 819 -1149 853
rect -1063 819 -1047 853
rect -1007 819 -991 853
rect -905 819 -889 853
rect -849 819 -833 853
rect -747 819 -731 853
rect -691 819 -675 853
rect -589 819 -573 853
rect -533 819 -517 853
rect -431 819 -415 853
rect -375 819 -359 853
rect -273 819 -257 853
rect -217 819 -201 853
rect -115 819 -99 853
rect -59 819 -43 853
rect 43 819 59 853
rect 99 819 115 853
rect 201 819 217 853
rect 257 819 273 853
rect 359 819 375 853
rect 415 819 431 853
rect 517 819 533 853
rect 573 819 589 853
rect 675 819 691 853
rect 731 819 747 853
rect 833 819 849 853
rect 889 819 905 853
rect 991 819 1007 853
rect 1047 819 1063 853
rect 1149 819 1165 853
rect 1205 819 1221 853
rect 1307 819 1323 853
rect 1363 819 1379 853
rect 1465 819 1481 853
rect 1521 819 1537 853
rect -1922 478 -1762 700
rect 1762 478 1922 700
rect -2322 118 -2162 340
rect 2162 118 2322 340
rect -2322 -940 -2162 -718
rect 2162 -940 2322 -718
rect -1922 -1300 -1762 -1078
rect 1762 -1300 1922 -1078
rect -1537 -1462 -1521 -1428
rect -1481 -1462 -1465 -1428
rect -1379 -1462 -1363 -1428
rect -1323 -1462 -1307 -1428
rect -1221 -1462 -1205 -1428
rect -1165 -1462 -1149 -1428
rect -1063 -1462 -1047 -1428
rect -1007 -1462 -991 -1428
rect -905 -1462 -889 -1428
rect -849 -1462 -833 -1428
rect -747 -1462 -731 -1428
rect -691 -1462 -675 -1428
rect -589 -1462 -573 -1428
rect -533 -1462 -517 -1428
rect -431 -1462 -415 -1428
rect -375 -1462 -359 -1428
rect -273 -1462 -257 -1428
rect -217 -1462 -201 -1428
rect -115 -1462 -99 -1428
rect -59 -1462 -43 -1428
rect 43 -1462 59 -1428
rect 99 -1462 115 -1428
rect 201 -1462 217 -1428
rect 257 -1462 273 -1428
rect 359 -1462 375 -1428
rect 415 -1462 431 -1428
rect 517 -1462 533 -1428
rect 573 -1462 589 -1428
rect 675 -1462 691 -1428
rect 731 -1462 747 -1428
rect 833 -1462 849 -1428
rect 889 -1462 905 -1428
rect 991 -1462 1007 -1428
rect 1047 -1462 1063 -1428
rect 1149 -1462 1165 -1428
rect 1205 -1462 1221 -1428
rect 1307 -1462 1323 -1428
rect 1363 -1462 1379 -1428
rect 1465 -1462 1481 -1428
rect 1521 -1462 1537 -1428
rect -1597 -1512 -1563 -1496
rect -1597 -2504 -1563 -2488
rect -1439 -1512 -1405 -1496
rect -1439 -2504 -1405 -2488
rect -1281 -1512 -1247 -1496
rect -1281 -2504 -1247 -2488
rect -1123 -1512 -1089 -1496
rect -1123 -2504 -1089 -2488
rect -965 -1512 -931 -1496
rect -965 -2504 -931 -2488
rect -807 -1512 -773 -1496
rect -807 -2504 -773 -2488
rect -649 -1512 -615 -1496
rect -649 -2504 -615 -2488
rect -491 -1512 -457 -1496
rect -491 -2504 -457 -2488
rect -333 -1512 -299 -1496
rect -333 -2504 -299 -2488
rect -175 -1512 -141 -1496
rect -175 -2504 -141 -2488
rect -17 -1512 17 -1496
rect -17 -2504 17 -2488
rect 141 -1512 175 -1496
rect 141 -2504 175 -2488
rect 299 -1512 333 -1496
rect 299 -2504 333 -2488
rect 457 -1512 491 -1496
rect 457 -2504 491 -2488
rect 615 -1512 649 -1496
rect 615 -2504 649 -2488
rect 773 -1512 807 -1496
rect 773 -2504 807 -2488
rect 931 -1512 965 -1496
rect 931 -2504 965 -2488
rect 1089 -1512 1123 -1496
rect 1089 -2504 1123 -2488
rect 1247 -1512 1281 -1496
rect 1247 -2504 1281 -2488
rect 1405 -1512 1439 -1496
rect 1405 -2504 1439 -2488
rect 1563 -1512 1597 -1496
rect 1563 -2504 1597 -2488
rect -1922 -2922 -1762 -2700
rect 1762 -2922 1922 -2700
rect -2322 -3322 -2162 -3100
rect 2162 -3322 2322 -3100
<< viali >>
rect -2162 2562 -2100 2722
rect -2100 2562 2100 2722
rect 2100 2562 2162 2722
rect -2322 392 -2162 2448
rect -1762 2162 -1700 2322
rect -1700 2162 1700 2322
rect 1700 2162 1762 2322
rect -1922 714 -1762 2086
rect -1603 1947 -1521 1981
rect -1521 1947 -1481 1981
rect -1481 1947 -1363 1981
rect -1363 1947 -1323 1981
rect -1323 1947 -1205 1981
rect -1205 1947 -1165 1981
rect -1165 1947 -1047 1981
rect -1047 1947 -1007 1981
rect -1007 1947 -889 1981
rect -889 1947 -849 1981
rect -849 1947 -731 1981
rect -731 1947 -691 1981
rect -691 1947 -573 1981
rect -573 1947 -533 1981
rect -533 1947 -415 1981
rect -415 1947 -375 1981
rect -375 1947 -257 1981
rect -257 1947 -217 1981
rect -217 1947 -99 1981
rect -99 1947 -59 1981
rect -59 1947 59 1981
rect 59 1947 99 1981
rect 99 1947 217 1981
rect 217 1947 257 1981
rect 257 1947 375 1981
rect 375 1947 415 1981
rect 415 1947 533 1981
rect 533 1947 573 1981
rect 573 1947 691 1981
rect 691 1947 731 1981
rect 731 1947 849 1981
rect 849 1947 889 1981
rect 889 1947 1007 1981
rect 1007 1947 1047 1981
rect 1047 1947 1165 1981
rect 1165 1947 1205 1981
rect 1205 1947 1323 1981
rect 1323 1947 1363 1981
rect 1363 1947 1481 1981
rect 1481 1947 1521 1981
rect 1521 1947 1603 1981
rect -1597 912 -1563 1888
rect -1439 912 -1405 1888
rect -1281 912 -1247 1888
rect -1123 912 -1089 1888
rect -965 912 -931 1888
rect -807 912 -773 1888
rect -649 912 -615 1888
rect -491 912 -457 1888
rect -333 912 -299 1888
rect -175 912 -141 1888
rect -17 912 17 1888
rect 141 912 175 1888
rect 299 912 333 1888
rect 457 912 491 1888
rect 615 912 649 1888
rect 773 912 807 1888
rect 931 912 965 1888
rect 1089 912 1123 1888
rect 1247 912 1281 1888
rect 1405 912 1439 1888
rect 1563 912 1597 1888
rect 1762 714 1922 2086
rect -1762 478 -1700 638
rect -1700 478 1700 638
rect 1700 478 1762 638
rect 2162 392 2322 2448
rect -2162 118 -2100 278
rect -2100 118 2100 278
rect 2100 118 2162 278
rect -2162 -878 -2100 -718
rect -2100 -878 2100 -718
rect 2100 -878 2162 -718
rect -2322 -3048 -2162 -992
rect -1762 -1238 -1700 -1078
rect -1700 -1238 1700 -1078
rect 1700 -1238 1762 -1078
rect -1922 -2686 -1762 -1314
rect -1597 -2488 -1563 -1512
rect -1439 -2488 -1405 -1512
rect -1281 -2488 -1247 -1512
rect -1123 -2488 -1089 -1512
rect -965 -2488 -931 -1512
rect -807 -2488 -773 -1512
rect -649 -2488 -615 -1512
rect -491 -2488 -457 -1512
rect -333 -2488 -299 -1512
rect -175 -2488 -141 -1512
rect -17 -2488 17 -1512
rect 141 -2488 175 -1512
rect 299 -2488 333 -1512
rect 457 -2488 491 -1512
rect 615 -2488 649 -1512
rect 773 -2488 807 -1512
rect 931 -2488 965 -1512
rect 1089 -2488 1123 -1512
rect 1247 -2488 1281 -1512
rect 1405 -2488 1439 -1512
rect 1563 -2488 1597 -1512
rect -1603 -2572 -1521 -2538
rect -1521 -2572 -1481 -2538
rect -1481 -2572 -1363 -2538
rect -1363 -2572 -1323 -2538
rect -1323 -2572 -1205 -2538
rect -1205 -2572 -1165 -2538
rect -1165 -2572 -1047 -2538
rect -1047 -2572 -1007 -2538
rect -1007 -2572 -889 -2538
rect -889 -2572 -849 -2538
rect -849 -2572 -731 -2538
rect -731 -2572 -691 -2538
rect -691 -2572 -573 -2538
rect -573 -2572 -533 -2538
rect -533 -2572 -415 -2538
rect -415 -2572 -375 -2538
rect -375 -2572 -257 -2538
rect -257 -2572 -217 -2538
rect -217 -2572 -99 -2538
rect -99 -2572 -59 -2538
rect -59 -2572 59 -2538
rect 59 -2572 99 -2538
rect 99 -2572 217 -2538
rect 217 -2572 257 -2538
rect 257 -2572 375 -2538
rect 375 -2572 415 -2538
rect 415 -2572 533 -2538
rect 533 -2572 573 -2538
rect 573 -2572 691 -2538
rect 691 -2572 731 -2538
rect 731 -2572 849 -2538
rect 849 -2572 889 -2538
rect 889 -2572 1007 -2538
rect 1007 -2572 1047 -2538
rect 1047 -2572 1165 -2538
rect 1165 -2572 1205 -2538
rect 1205 -2572 1323 -2538
rect 1323 -2572 1363 -2538
rect 1363 -2572 1481 -2538
rect 1481 -2572 1521 -2538
rect 1521 -2572 1603 -2538
rect 1762 -2686 1922 -1314
rect -1762 -2922 -1700 -2762
rect -1700 -2922 1700 -2762
rect 1700 -2922 1762 -2762
rect 2162 -3048 2322 -992
rect -2162 -3322 -2100 -3162
rect -2100 -3322 2100 -3162
rect 2100 -3322 2162 -3162
<< metal1 >>
rect -2328 2722 2328 2728
rect -2328 2562 -2162 2722
rect 2162 2562 2328 2722
rect -2328 2460 2328 2562
rect -2328 2448 -2060 2460
rect -2328 392 -2322 2448
rect -2162 392 -2060 2448
rect 2060 2448 2328 2460
rect -2001 2340 2000 2400
rect -2001 2119 -1941 2340
rect 1940 2119 2000 2340
rect -2001 2086 2000 2119
rect -2001 2059 -1922 2086
rect -2000 714 -1922 2059
rect -1762 2059 1762 2086
rect -1762 734 -1660 2059
rect -1603 1987 -1557 2059
rect -1287 1987 -1241 2059
rect -971 1987 -925 2059
rect -655 1987 -609 2059
rect -339 1987 -293 2059
rect -23 1987 23 2059
rect 293 1987 339 2059
rect 609 1987 655 2059
rect 925 1987 971 2059
rect 1241 1987 1287 2059
rect 1557 1987 1603 2059
rect -1615 1981 1615 1987
rect -1615 1947 -1603 1981
rect 1603 1947 1615 1981
rect -1615 1941 1615 1947
rect -1603 1888 -1557 1941
rect -1603 912 -1597 1888
rect -1563 912 -1557 1888
rect -1603 900 -1557 912
rect -1445 1888 -1399 1900
rect -1445 912 -1439 1888
rect -1405 912 -1399 1888
rect -1445 864 -1399 912
rect -1287 1888 -1241 1941
rect -1287 912 -1281 1888
rect -1247 912 -1241 1888
rect -1287 900 -1241 912
rect -1129 1888 -1083 1900
rect -1129 912 -1123 1888
rect -1089 912 -1083 1888
rect -1129 864 -1083 912
rect -971 1888 -925 1941
rect -971 912 -965 1888
rect -931 912 -925 1888
rect -971 900 -925 912
rect -813 1888 -767 1900
rect -813 912 -807 1888
rect -773 912 -767 1888
rect -813 864 -767 912
rect -655 1888 -609 1941
rect -655 912 -649 1888
rect -615 912 -609 1888
rect -655 900 -609 912
rect -497 1888 -451 1900
rect -497 912 -491 1888
rect -457 912 -451 1888
rect -497 864 -451 912
rect -339 1888 -293 1941
rect -339 912 -333 1888
rect -299 912 -293 1888
rect -339 900 -293 912
rect -181 1888 -135 1900
rect -181 912 -175 1888
rect -141 912 -135 1888
rect -181 864 -135 912
rect -23 1888 23 1941
rect -23 912 -17 1888
rect 17 912 23 1888
rect -23 900 23 912
rect 135 1888 181 1900
rect 135 912 141 1888
rect 175 912 181 1888
rect 135 864 181 912
rect 293 1888 339 1941
rect 293 912 299 1888
rect 333 912 339 1888
rect 293 900 339 912
rect 451 1888 497 1900
rect 451 912 457 1888
rect 491 912 497 1888
rect 451 864 497 912
rect 609 1888 655 1941
rect 609 912 615 1888
rect 649 912 655 1888
rect 609 900 655 912
rect 767 1888 813 1900
rect 767 912 773 1888
rect 807 912 813 1888
rect 767 864 813 912
rect 925 1888 971 1941
rect 925 912 931 1888
rect 965 912 971 1888
rect 925 900 971 912
rect 1083 1888 1129 1900
rect 1083 912 1089 1888
rect 1123 912 1129 1888
rect 1083 864 1129 912
rect 1241 1888 1287 1941
rect 1241 912 1247 1888
rect 1281 912 1287 1888
rect 1241 900 1287 912
rect 1399 1888 1445 1900
rect 1399 912 1405 1888
rect 1439 912 1445 1888
rect 1399 864 1445 912
rect 1557 1888 1603 1941
rect 1557 912 1563 1888
rect 1597 912 1603 1888
rect 1557 900 1603 912
rect -1445 858 1445 864
rect -1449 780 -1439 858
rect 1439 780 1449 858
rect -1445 774 1445 780
rect 1650 734 1762 2059
rect -1762 714 1762 734
rect 1922 714 2000 2086
rect -2000 638 2000 714
rect -2000 478 -1762 638
rect 1762 478 2000 638
rect -2000 400 2000 478
rect -2328 340 -2060 392
rect 2060 392 2162 2448
rect 2322 392 2328 2448
rect 2060 340 2328 392
rect -2328 278 2328 340
rect -2328 118 -2162 278
rect 2162 118 2328 278
rect -2328 -718 2328 118
rect -2328 -878 -2162 -718
rect 2162 -878 2328 -718
rect -2328 -992 2328 -878
rect -2328 -2814 -2322 -992
rect -2162 -1078 2162 -992
rect -2162 -1238 -1762 -1078
rect 1762 -1238 2162 -1078
rect -2162 -1244 2162 -1238
rect -2162 -1314 -1756 -1244
rect -2162 -2686 -1922 -1314
rect -1762 -2686 -1756 -1314
rect -1445 -1316 1445 -1310
rect 1756 -1314 2162 -1244
rect -1449 -1394 -1439 -1316
rect 1439 -1394 1449 -1316
rect -1445 -1400 1445 -1394
rect -1603 -1512 -1557 -1500
rect -1603 -2488 -1597 -1512
rect -1563 -2488 -1557 -1512
rect -1603 -2532 -1557 -2488
rect -1445 -1512 -1399 -1400
rect -1445 -2488 -1439 -1512
rect -1405 -2488 -1399 -1512
rect -1445 -2500 -1399 -2488
rect -1287 -1512 -1241 -1500
rect -1287 -2488 -1281 -1512
rect -1247 -2488 -1241 -1512
rect -1287 -2532 -1241 -2488
rect -1129 -1512 -1083 -1400
rect -1129 -2488 -1123 -1512
rect -1089 -2488 -1083 -1512
rect -1129 -2500 -1083 -2488
rect -971 -1512 -925 -1500
rect -971 -2488 -965 -1512
rect -931 -2488 -925 -1512
rect -971 -2532 -925 -2488
rect -813 -1512 -767 -1400
rect -813 -2488 -807 -1512
rect -773 -2488 -767 -1512
rect -813 -2500 -767 -2488
rect -655 -1512 -609 -1500
rect -655 -2488 -649 -1512
rect -615 -2488 -609 -1512
rect -655 -2532 -609 -2488
rect -497 -1512 -451 -1400
rect -497 -2488 -491 -1512
rect -457 -2488 -451 -1512
rect -497 -2500 -451 -2488
rect -339 -1512 -293 -1500
rect -339 -2488 -333 -1512
rect -299 -2488 -293 -1512
rect -339 -2532 -293 -2488
rect -181 -1512 -135 -1400
rect -181 -2488 -175 -1512
rect -141 -2488 -135 -1512
rect -181 -2500 -135 -2488
rect -23 -1512 23 -1500
rect -23 -2488 -17 -1512
rect 17 -2488 23 -1512
rect -23 -2532 23 -2488
rect 135 -1512 181 -1400
rect 135 -2488 141 -1512
rect 175 -2488 181 -1512
rect 135 -2500 181 -2488
rect 293 -1512 339 -1500
rect 293 -2488 299 -1512
rect 333 -2488 339 -1512
rect 293 -2532 339 -2488
rect 451 -1512 497 -1400
rect 451 -2488 457 -1512
rect 491 -2488 497 -1512
rect 451 -2500 497 -2488
rect 609 -1512 655 -1500
rect 609 -2488 615 -1512
rect 649 -2488 655 -1512
rect 609 -2532 655 -2488
rect 767 -1512 813 -1400
rect 767 -2488 773 -1512
rect 807 -2488 813 -1512
rect 767 -2500 813 -2488
rect 925 -1512 971 -1500
rect 925 -2488 931 -1512
rect 965 -2488 971 -1512
rect 925 -2532 971 -2488
rect 1083 -1512 1129 -1400
rect 1083 -2488 1089 -1512
rect 1123 -2488 1129 -1512
rect 1083 -2500 1129 -2488
rect 1241 -1512 1287 -1500
rect 1241 -2488 1247 -1512
rect 1281 -2488 1287 -1512
rect 1241 -2532 1287 -2488
rect 1399 -1512 1445 -1400
rect 1399 -2488 1405 -1512
rect 1439 -2488 1445 -1512
rect 1399 -2500 1445 -2488
rect 1557 -1512 1603 -1500
rect 1557 -2488 1563 -1512
rect 1597 -2488 1603 -1512
rect 1557 -2532 1603 -2488
rect -1615 -2538 1615 -2532
rect -1615 -2572 -1603 -2538
rect 1603 -2572 1615 -2538
rect -1615 -2578 1615 -2572
rect -2162 -2755 -1756 -2686
rect -1603 -2755 -1557 -2578
rect -1287 -2755 -1241 -2578
rect -971 -2755 -925 -2578
rect -655 -2755 -609 -2578
rect -339 -2755 -293 -2578
rect -23 -2755 23 -2578
rect 293 -2755 339 -2578
rect 609 -2755 655 -2578
rect 925 -2755 971 -2578
rect 1241 -2755 1287 -2578
rect 1557 -2755 1603 -2578
rect 1756 -2686 1762 -1314
rect 1922 -2686 2162 -1314
rect 1756 -2755 2162 -2686
rect -2162 -2762 2162 -2755
rect -2162 -2814 -1762 -2762
rect 1762 -2814 2162 -2762
rect 2322 -2814 2328 -992
rect -2350 -3340 -2340 -2814
rect 2340 -3340 2350 -2814
<< via1 >>
rect -1941 2322 1940 2340
rect -1941 2162 -1762 2322
rect -1762 2162 1762 2322
rect 1762 2162 1940 2322
rect -1941 2119 1940 2162
rect -1439 780 1439 858
rect -1439 -1394 1439 -1316
rect -2340 -3048 -2322 -2814
rect -2322 -3048 -2162 -2814
rect -2162 -2922 -1762 -2814
rect -1762 -2922 1762 -2814
rect 1762 -2922 2162 -2814
rect -2162 -3048 2162 -2922
rect 2162 -3048 2322 -2814
rect 2322 -3048 2340 -2814
rect -2340 -3162 2340 -3048
rect -2340 -3322 -2162 -3162
rect -2162 -3322 2162 -3162
rect 2162 -3322 2340 -3162
rect -2340 -3340 2340 -3322
<< metal2 >>
rect -2400 2340 2400 2800
rect -2400 2119 -1941 2340
rect 1940 2119 2400 2340
rect -2400 2000 2400 2119
rect -1439 858 1439 868
rect -1439 -100 1439 780
rect -2400 -500 2400 -100
rect -1439 -1316 1439 -500
rect -1439 -1404 1439 -1394
rect -2400 -2814 2400 -2600
rect -2400 -3340 -2340 -2814
rect 2340 -3340 2400 -2814
rect -2400 -3400 2400 -3340
<< labels >>
flabel metal2 -2400 2000 -2395 2800 3 FreeSans 400 0 0 0 vdd
port 2 e
flabel metal2 -2400 -3400 -2395 -2600 3 FreeSans 400 0 0 0 vss
port 3 e
flabel metal2 -2400 -500 -2395 -100 3 FreeSans 400 0 0 0 clamp
port 1 e
<< end >>
