magic
tech sky130A
magscale 1 2
timestamp 1623205543
<< metal1 >>
rect -20400 3360 20500 49600
rect -199 505 201 565
rect -199 441 -139 505
rect -200 225 -139 441
rect 141 225 201 505
rect -200 165 201 225
rect -200 41 200 165
rect -206 -1632 -200 -1232
rect 200 -1632 206 -1232
rect -85199 -30024 -23576 -9757
rect -21510 -29400 -21500 -13300
rect -21160 -29400 -21150 -13300
rect -15450 -29400 -15440 -13300
rect -15100 -29400 -15090 -13300
rect 14490 -29400 14500 -13300
rect 14840 -29400 14850 -13300
rect 20550 -29400 20560 -13300
rect 20900 -29400 20910 -13300
rect -85209 -32280 -85199 -30024
rect -23576 -32280 -23566 -30024
<< via1 >>
rect -139 225 141 505
rect -200 -1632 200 -1232
rect -21500 -29400 -21160 -13300
rect -15440 -29400 -15100 -13300
rect 14500 -29400 14840 -13300
rect 20560 -29400 20900 -13300
rect -85199 -32280 -23576 -30024
<< metal2 >>
rect -20400 3360 20500 49600
rect 67695 40505 68695 40515
rect 67695 39495 68695 39505
rect 67695 36505 68695 36515
rect 67695 35495 68695 35505
rect 67695 32505 68695 32515
rect 67695 31495 68695 31505
rect 67695 28505 68695 28515
rect 67695 27495 68695 27505
rect 67695 24505 68695 24515
rect 67695 23495 68695 23505
rect 67695 20505 68695 20515
rect 67695 19495 68695 19505
rect 67695 16505 68695 16515
rect 67695 15495 68695 15505
rect 67695 12505 68695 12515
rect 67695 11495 68695 11505
rect 67695 8505 68695 8515
rect 67695 7495 68695 7505
rect 67695 4505 68695 4515
rect 67695 3495 68695 3505
rect -20400 2226 -4599 2426
rect -20400 1722 -20200 2226
rect -19456 1722 -4599 2226
rect -20400 1522 -4599 1722
rect -6553 1422 -6453 1522
rect -22348 422 -16669 423
rect -22350 -50 -16669 422
rect -22822 -1386 -16669 -50
rect -22342 -1388 -16669 -1386
rect -85199 -30024 -23576 -9757
rect -21900 -13290 -21160 -13280
rect -18340 -13418 -16669 -1388
rect -15440 -13300 -14700 -13290
rect -21900 -29420 -21160 -29410
rect -16566 -29414 -16506 -28852
rect -85199 -32290 -23576 -32280
rect -16682 -29474 -16506 -29414
rect -16462 -29415 -16402 -28852
rect -15440 -29410 -14700 -29400
rect -16682 -64204 -16622 -29474
rect -16462 -29475 -16262 -29415
rect -16322 -64204 -16262 -29475
rect -6553 -64204 -6453 1322
rect -5503 -64204 -4599 1522
rect -139 505 141 515
rect -139 215 141 225
rect -200 -1232 200 -1226
rect -3100 -4600 -2300 -4590
rect -200 -5000 200 -1632
rect 2300 -4600 3100 -4590
rect -3100 -9410 -2300 -9400
rect -200 -64204 200 -9000
rect 3539 -5133 15510 3360
rect 67695 505 68695 515
rect 3539 -5543 15510 -5533
rect 17660 -377 22100 422
rect 17660 -1267 22922 -377
rect 67695 -505 68695 -495
rect 2300 -9410 3100 -9400
rect 14100 -13290 14840 -13280
rect 17660 -13400 19331 -1267
rect 67695 -3495 68695 -3485
rect 67695 -4505 68695 -4495
rect 25693 -5497 26693 -5487
rect 25693 -6507 26693 -6497
rect 29695 -5495 30695 -5485
rect 29695 -6505 30695 -6495
rect 33695 -5495 34695 -5485
rect 33695 -6505 34695 -6495
rect 37695 -5495 38695 -5485
rect 37695 -6505 38695 -6495
rect 41695 -5495 42695 -5485
rect 41695 -6505 42695 -6495
rect 45695 -5495 46695 -5485
rect 45695 -6505 46695 -6495
rect 49695 -5495 50695 -5485
rect 49695 -6505 50695 -6495
rect 53695 -5495 54695 -5485
rect 53695 -6505 54695 -6495
rect 57695 -5495 58695 -5485
rect 57695 -6505 58695 -6495
rect 61695 -5495 62695 -5485
rect 61695 -6505 62695 -6495
rect 65695 -5495 66695 -5485
rect 65695 -6505 66695 -6495
rect 20560 -13300 21300 -13290
rect 19434 -28994 19494 -28852
rect 14100 -29420 14840 -29410
rect 19317 -29054 19494 -28994
rect 19538 -28999 19598 -28852
rect 19317 -64204 19377 -29054
rect 19538 -29059 19797 -28999
rect 19737 -64204 19797 -29059
rect 20560 -29410 21300 -29400
<< rmetal2 >>
rect -6553 1322 -6453 1422
<< via2 >>
rect 67695 39505 68695 40505
rect 67695 35505 68695 36505
rect 67695 31505 68695 32505
rect 67695 27505 68695 28505
rect 67695 23505 68695 24505
rect 67695 19505 68695 20505
rect 67695 15505 68695 16505
rect 67695 11505 68695 12505
rect 67695 7505 68695 8505
rect 67695 3505 68695 4505
rect -20200 1722 -19456 2226
rect -21900 -13300 -21160 -13290
rect -21900 -29400 -21500 -13300
rect -21500 -29400 -21160 -13300
rect -21900 -29410 -21160 -29400
rect -85199 -32280 -23576 -30024
rect -15440 -29400 -15100 -13300
rect -15100 -29400 -14700 -13300
rect -139 225 141 505
rect -3100 -9400 -2300 -4600
rect 2300 -9400 3100 -4600
rect 3539 -5533 15510 -5133
rect 67695 -495 68695 505
rect 14100 -13300 14840 -13290
rect 14100 -29400 14500 -13300
rect 14500 -29400 14840 -13300
rect 67695 -4495 68695 -3495
rect 25693 -6497 26693 -5497
rect 29695 -6495 30695 -5495
rect 33695 -6495 34695 -5495
rect 37695 -6495 38695 -5495
rect 41695 -6495 42695 -5495
rect 45695 -6495 46695 -5495
rect 49695 -6495 50695 -5495
rect 53695 -6495 54695 -5495
rect 57695 -6495 58695 -5495
rect 61695 -6495 62695 -5495
rect 65695 -6495 66695 -5495
rect 14100 -29410 14840 -29400
rect 20560 -29400 20900 -13300
rect 20900 -29400 21300 -13300
<< metal3 >>
rect -119200 -4000 -79200 66802
rect -75200 56800 62100 66800
rect -18400 43600 62100 56800
rect -18400 3300 18500 43600
rect 64100 40505 96100 41200
rect 64100 39600 67695 40505
rect 66100 39505 67695 39600
rect 68695 39505 96100 40505
rect 66100 36505 96100 39505
rect 66100 35505 67695 36505
rect 68695 35505 96100 36505
rect 66100 32505 96100 35505
rect 66100 31505 67695 32505
rect 68695 31505 96100 32505
rect 66100 28505 96100 31505
rect 66100 27505 67695 28505
rect 68695 27505 96100 28505
rect 66100 24505 96100 27505
rect 66100 23505 67695 24505
rect 68695 23505 96100 24505
rect 66100 20505 96100 23505
rect 66100 19505 67695 20505
rect 68695 19505 96100 20505
rect 66100 16505 96100 19505
rect 66100 15505 67695 16505
rect 68695 15505 96100 16505
rect 66100 12505 96100 15505
rect 66100 11505 67695 12505
rect 68695 11505 96100 12505
rect 66100 8505 96100 11505
rect 66100 7505 67695 8505
rect 68695 7505 96100 8505
rect 66100 4505 96100 7505
rect -20400 2226 -19256 2426
rect -20400 1722 -20200 2226
rect -19456 1722 -19256 2226
rect -20400 1522 -19256 1722
rect -200 505 202 3300
rect 18501 1522 20501 3519
rect 66100 3505 67695 4505
rect 68695 3505 96100 4505
rect -200 225 -139 505
rect 141 225 202 505
rect -200 162 202 225
rect 66100 505 96100 3505
rect 66100 -495 67695 505
rect 68695 -495 96100 505
rect 2278 -4000 22640 -2000
rect 66100 -3495 96100 -495
rect 66100 -4000 67695 -3495
rect -119200 -4576 -22388 -4000
rect 2278 -4495 67695 -4000
rect 68695 -4495 96100 -3495
rect 2278 -4576 96100 -4495
rect -119200 -4600 -2276 -4576
rect -119200 -9400 -3100 -4600
rect -2300 -9400 -2276 -4600
rect -119200 -11348 -2276 -9400
rect 2276 -4600 96100 -4576
rect 2276 -9400 2300 -4600
rect 3100 -5133 96100 -4600
rect 3100 -5533 3539 -5133
rect 15510 -5495 96100 -5133
rect 15510 -5497 29695 -5495
rect 15510 -5533 25693 -5497
rect 3100 -6497 25693 -5533
rect 26693 -6495 29695 -5497
rect 30695 -6495 33695 -5495
rect 34695 -6495 37695 -5495
rect 38695 -6495 41695 -5495
rect 42695 -6495 45695 -5495
rect 46695 -6495 49695 -5495
rect 50695 -6495 53695 -5495
rect 54695 -6495 57695 -5495
rect 58695 -6495 61695 -5495
rect 62695 -6495 65695 -5495
rect 66695 -6495 96100 -5495
rect 26693 -6497 96100 -6495
rect 3100 -9400 96100 -6497
rect 2276 -9424 96100 -9400
rect -119200 -13290 -21135 -11348
rect -7924 -13266 -2276 -11348
rect 2278 -11647 96100 -9424
rect -119200 -24000 -21900 -13290
rect -22443 -29410 -21900 -24000
rect -21160 -29410 -21135 -13290
rect -22443 -29433 -21135 -29410
rect -15464 -13300 -11464 -13276
rect -15464 -29400 -15440 -13300
rect -14700 -29400 -11464 -13300
rect -85209 -30024 -23566 -30019
rect -15464 -30024 -11464 -29400
rect -7924 -13290 14864 -13266
rect 22500 -13276 96100 -11647
rect -7924 -29410 14100 -13290
rect 14840 -29410 14864 -13290
rect 21164 -13295 96100 -13276
rect 20550 -13300 96100 -13295
rect 20550 -29400 20560 -13300
rect 21300 -29400 96100 -13300
rect 20550 -29405 96100 -29400
rect -7924 -29434 14864 -29410
rect 21164 -29424 96100 -29405
rect 22500 -30024 96100 -29424
rect -119200 -32280 -85199 -30024
rect -23576 -32280 96100 -30024
rect -119200 -64000 96100 -32280
<< via3 >>
rect 67695 39505 68695 40505
rect 67695 35505 68695 36505
rect 67695 31505 68695 32505
rect 67695 27505 68695 28505
rect 67695 23505 68695 24505
rect 67695 19505 68695 20505
rect 67695 15505 68695 16505
rect 67695 11505 68695 12505
rect 67695 7505 68695 8505
rect -20200 1722 -19456 2226
rect 67695 3505 68695 4505
rect -139 225 141 505
rect 67695 -495 68695 505
rect 67695 -4495 68695 -3495
rect -3100 -9400 -2300 -4600
rect 2300 -9400 3100 -4600
rect 3539 -5533 15510 -5133
rect 25693 -6497 26693 -5497
rect 29695 -6495 30695 -5495
rect 33695 -6495 34695 -5495
rect 37695 -6495 38695 -5495
rect 41695 -6495 42695 -5495
rect 45695 -6495 46695 -5495
rect 49695 -6495 50695 -5495
rect 53695 -6495 54695 -5495
rect 57695 -6495 58695 -5495
rect 61695 -6495 62695 -5495
rect 65695 -6495 66695 -5495
rect -21900 -29410 -21160 -13290
rect -15440 -29400 -14700 -13300
rect 14100 -29410 14840 -13290
rect 20560 -29400 21300 -13300
rect -85199 -32280 -23576 -30024
<< metal4 >>
rect -119200 -4000 -79200 66802
rect -75200 56800 62100 66800
rect -18400 43600 62100 56800
rect -18400 3300 18500 43600
rect 64100 40505 96100 41200
rect 64100 39600 67695 40505
rect 66100 39505 67695 39600
rect 68695 39505 96100 40505
rect 66100 36505 96100 39505
rect 66100 35505 67695 36505
rect 68695 35505 96100 36505
rect 66100 32505 96100 35505
rect 66100 31505 67695 32505
rect 68695 31505 96100 32505
rect 66100 28505 96100 31505
rect 66100 27505 67695 28505
rect 68695 27505 96100 28505
rect 66100 24505 96100 27505
rect 66100 23505 67695 24505
rect 68695 23505 96100 24505
rect 66100 20505 96100 23505
rect 66100 19505 67695 20505
rect 68695 19505 96100 20505
rect 66100 16505 96100 19505
rect 66100 15505 67695 16505
rect 68695 15505 96100 16505
rect 66100 12505 96100 15505
rect 66100 11505 67695 12505
rect 68695 11505 96100 12505
rect 66100 8505 96100 11505
rect 66100 7505 67695 8505
rect 68695 7505 96100 8505
rect 66100 4505 96100 7505
rect -20400 2256 -19256 2426
rect -20400 1834 -20300 2256
rect -19356 1834 -19256 2256
rect -20400 1722 -20200 1834
rect -19456 1722 -19256 1834
rect -20400 1522 -19256 1722
rect -200 505 202 3300
rect 18501 1522 20501 3519
rect 66100 3505 67695 4505
rect 68695 3505 96100 4505
rect -200 225 -139 505
rect 141 225 202 505
rect -200 162 202 225
rect 66100 505 96100 3505
rect 66100 -495 67695 505
rect 68695 -495 96100 505
rect 2278 -4000 22640 -2000
rect 66100 -3495 96100 -495
rect 66100 -4000 67695 -3495
rect -119200 -4576 -22388 -4000
rect 2278 -4495 67695 -4000
rect 68695 -4495 96100 -3495
rect 2278 -4576 96100 -4495
rect -119200 -4600 -2276 -4576
rect -119200 -9400 -3100 -4600
rect -2300 -9400 -2276 -4600
rect -119200 -11348 -2276 -9400
rect 2276 -4600 96100 -4576
rect 2276 -9400 2300 -4600
rect 3100 -5133 96100 -4600
rect 3100 -5533 3539 -5133
rect 15510 -5495 96100 -5133
rect 15510 -5497 29695 -5495
rect 15510 -5533 25693 -5497
rect 3100 -6497 25693 -5533
rect 26693 -6495 29695 -5497
rect 30695 -6495 33695 -5495
rect 34695 -6495 37695 -5495
rect 38695 -6495 41695 -5495
rect 42695 -6495 45695 -5495
rect 46695 -6495 49695 -5495
rect 50695 -6495 53695 -5495
rect 54695 -6495 57695 -5495
rect 58695 -6495 61695 -5495
rect 62695 -6495 65695 -5495
rect 66695 -6495 96100 -5495
rect 26693 -6497 96100 -6495
rect 3100 -9400 96100 -6497
rect 2276 -9424 96100 -9400
rect -119200 -13290 -21135 -11348
rect -7924 -13266 -2276 -11348
rect 2278 -11647 96100 -9424
rect -119200 -24000 -21900 -13290
rect -22443 -29410 -21900 -24000
rect -21160 -29410 -21135 -13290
rect -22443 -29433 -21135 -29410
rect -15464 -13300 -11464 -13276
rect -15464 -29400 -15440 -13300
rect -14700 -29400 -11464 -13300
rect -85200 -30024 -23575 -30023
rect -15464 -30024 -11464 -29400
rect -7924 -13290 14864 -13266
rect 22500 -13276 96100 -11647
rect -7924 -29410 14100 -13290
rect 14840 -29410 14864 -13290
rect 21164 -13299 96100 -13276
rect 20559 -13300 96100 -13299
rect 20559 -29400 20560 -13300
rect 21300 -29400 96100 -13300
rect 20559 -29401 96100 -29400
rect -7924 -29434 14864 -29410
rect 21164 -29424 96100 -29401
rect 22500 -30024 96100 -29424
rect -119200 -32280 -85199 -30024
rect -23576 -32280 96100 -30024
rect -119200 -64000 96100 -32280
<< via4 >>
rect 67695 39505 68695 40505
rect 67695 35505 68695 36505
rect 67695 31505 68695 32505
rect 67695 27505 68695 28505
rect 67695 23505 68695 24505
rect 67695 19505 68695 20505
rect 67695 15505 68695 16505
rect 67695 11505 68695 12505
rect 67695 7505 68695 8505
rect -20300 2226 -19356 2256
rect -20300 1834 -20200 2226
rect -20200 1834 -19456 2226
rect -19456 1834 -19356 2226
rect 67695 3505 68695 4505
rect -139 225 141 505
rect 67695 -495 68695 505
rect 67695 -4495 68695 -3495
rect -3100 -9400 -2300 -4600
rect 2300 -9400 3100 -4600
rect 3539 -5533 15510 -5133
rect 25693 -6497 26693 -5497
rect 29695 -6495 30695 -5495
rect 33695 -6495 34695 -5495
rect 37695 -6495 38695 -5495
rect 41695 -6495 42695 -5495
rect 45695 -6495 46695 -5495
rect 49695 -6495 50695 -5495
rect 53695 -6495 54695 -5495
rect 57695 -6495 58695 -5495
rect 61695 -6495 62695 -5495
rect 65695 -6495 66695 -5495
rect -21900 -29410 -21160 -13290
rect -15440 -29400 -14700 -13300
rect 14100 -29410 14840 -13290
rect 20560 -29400 21300 -13300
rect -85199 -32280 -23576 -30024
<< metal5 >>
rect -119200 -4000 -79200 66802
rect -75200 56800 62100 66800
rect -18400 43600 62100 56800
rect -18400 3300 18500 43600
rect 64100 40505 96100 41200
rect 64100 39600 67695 40505
rect 66100 39505 67695 39600
rect 68695 39505 96100 40505
rect 66100 36505 96100 39505
rect 66100 35505 67695 36505
rect 68695 35505 96100 36505
rect 66100 32505 96100 35505
rect 66100 31505 67695 32505
rect 68695 31505 96100 32505
rect 66100 28505 96100 31505
rect 66100 27505 67695 28505
rect 68695 27505 96100 28505
rect 66100 24505 96100 27505
rect 66100 23505 67695 24505
rect 68695 23505 96100 24505
rect 66100 20505 96100 23505
rect 66100 19505 67695 20505
rect 68695 19505 96100 20505
rect 66100 16505 96100 19505
rect 66100 15505 67695 16505
rect 68695 15505 96100 16505
rect 66100 12505 96100 15505
rect 66100 11505 67695 12505
rect 68695 11505 96100 12505
rect 66100 8505 96100 11505
rect 66100 7505 67695 8505
rect 68695 7505 96100 8505
rect 66100 4505 96100 7505
rect -20400 2256 -19256 2356
rect -20400 1834 -20300 2256
rect -19356 1834 -19256 2256
rect -20400 1734 -19256 1834
rect -200 505 202 3300
rect 18501 1522 20501 3519
rect 66100 3505 67695 4505
rect 68695 3505 96100 4505
rect -200 225 -139 505
rect 141 225 202 505
rect -200 162 202 225
rect 66100 505 96100 3505
rect 66100 -495 67695 505
rect 68695 -495 96100 505
rect 2278 -4000 22640 -2000
rect 66100 -3495 96100 -495
rect 66100 -4000 67695 -3495
rect -119200 -4576 -22388 -4000
rect 2278 -4495 67695 -4000
rect 68695 -4495 96100 -3495
rect 2278 -4576 96100 -4495
rect -119200 -4600 -2276 -4576
rect -119200 -9400 -3100 -4600
rect -2300 -9400 -2276 -4600
rect -119200 -11348 -2276 -9400
rect 2276 -4600 96100 -4576
rect 2276 -9400 2300 -4600
rect 3100 -5133 96100 -4600
rect 3100 -5533 3539 -5133
rect 15510 -5495 96100 -5133
rect 15510 -5497 29695 -5495
rect 15510 -5533 25693 -5497
rect 3100 -6497 25693 -5533
rect 26693 -6495 29695 -5497
rect 30695 -6495 33695 -5495
rect 34695 -6495 37695 -5495
rect 38695 -6495 41695 -5495
rect 42695 -6495 45695 -5495
rect 46695 -6495 49695 -5495
rect 50695 -6495 53695 -5495
rect 54695 -6495 57695 -5495
rect 58695 -6495 61695 -5495
rect 62695 -6495 65695 -5495
rect 66695 -6495 96100 -5495
rect 26693 -6497 96100 -6495
rect 3100 -9400 96100 -6497
rect 2276 -9424 96100 -9400
rect -119200 -13290 -21135 -11348
rect -7924 -13266 -2276 -11348
rect 2278 -11647 96100 -9424
rect -119200 -24000 -21900 -13290
rect -22443 -29410 -21900 -24000
rect -21160 -29410 -21135 -13290
rect -22443 -29433 -21135 -29410
rect -15464 -13300 -11464 -13276
rect -15464 -29400 -15440 -13300
rect -14700 -29400 -11464 -13300
rect -21924 -29434 -21136 -29433
rect -85223 -30024 -23552 -30000
rect -15464 -30024 -11464 -29400
rect -7924 -13290 14864 -13266
rect 22500 -13276 96100 -11647
rect -7924 -29410 14100 -13290
rect 14840 -29410 14864 -13290
rect -7924 -29434 14864 -29410
rect 20536 -13300 96100 -13276
rect 20536 -29400 20560 -13300
rect 21300 -29400 96100 -13300
rect 20536 -29424 96100 -29400
rect 22500 -30024 96100 -29424
rect -119200 -32280 -85199 -30024
rect -23576 -32280 96100 -30024
rect -119200 -64000 96100 -32280
use sky130_fd_pr__res_generic_po_U6Z5S8  sky130_fd_pr__res_generic_po_U6Z5S8_0
timestamp 1623025674
transform 1 0 0 0 1 -600
box -200 -703 200 703
use nmos_waffle_36x36  nmos_waffle_36x36_0
timestamp 1622614837
transform 1 0 22500 0 1 0
box -10800 -10800 50400 50400
use pmos_waffle_48x48  pmos_waffle_48x48_0
timestamp 1622615317
transform -1 0 -22400 0 1 0
box -10800 -10800 63600 63600
use esd_cell_well  esd_cell_well_0
timestamp 1622610789
transform 0 -1 -300 1 0 -7000
box -2400 -3400 2400 2800
use gate_drive  gate_drive_0
timestamp 1621730769
transform 0 -1 -17500 1 0 -20900
box -8500 -2400 7600 4000
use gate_drive  gate_drive_1
timestamp 1621730769
transform 0 -1 18500 1 0 -20900
box -8500 -2400 7600 4000
<< labels >>
flabel metal2 -16682 -64204 -16622 -64203 1 FreeSans 400 0 0 0 p_in
port 3 n
flabel metal2 -16322 -64204 -16262 -64203 1 FreeSans 400 0 0 0 p_in_n
port 4 n
flabel metal2 -6553 -64204 -6453 -64202 1 FreeSans 400 0 0 0 ref_current_kelvin
port 6 n
flabel metal2 -5503 -64204 -4599 -64199 1 FreeSans 400 0 0 0 ref_current
port 5 n
flabel metal2 -200 -64204 200 -64199 1 FreeSans 400 0 0 0 sw_node_esd
port 8 n
flabel metal2 19317 -64204 19377 -64203 1 FreeSans 400 0 0 0 n_in
port 1 n
flabel metal2 19737 -64204 19797 -64203 1 FreeSans 400 0 0 0 n_in_n
port 2 n
flabel metal5 -75200 66764 62100 66800 1 FreeSans 8000 0 0 0 sw_node
port 7 n
flabel metal5 -119200 66800 -79200 66802 5 FreeSans 8000 0 0 0 vdd_pwr
port 9 s
flabel metal5 -119200 -64000 -119179 -30024 1 FreeSans 8000 0 0 0 vss
port 10 n
<< end >>
