magic
tech sky130A
magscale 1 2
timestamp 1623996740
<< nwell >>
rect -922 -5049 -826 -4529
rect 1000 -9000 11000 -4600
<< pwell >>
rect -992 -4435 -753 -4109
rect 1000 -4400 11000 0
<< mvpsubdiff >>
rect 1066 -78 10934 -66
rect 1066 -238 1300 -78
rect 10700 -238 10934 -78
rect 1066 -250 10934 -238
rect 1066 -300 1250 -250
rect 1066 -4100 1078 -300
rect 1238 -4100 1250 -300
rect -988 -4169 -760 -4135
rect 1066 -4150 1250 -4100
rect 10750 -300 10934 -250
rect 10750 -4100 10762 -300
rect 10922 -4100 10934 -300
rect 10750 -4150 10934 -4100
rect 1066 -4162 10934 -4150
rect 1066 -4322 1300 -4162
rect 10700 -4322 10934 -4162
rect 1066 -4334 10934 -4322
<< mvnsubdiff >>
rect 1066 -4678 10934 -4666
rect 1066 -4838 1300 -4678
rect 10700 -4838 10934 -4678
rect 1066 -4850 10934 -4838
rect 1066 -4900 1250 -4850
rect -988 -4983 -760 -4949
rect 1066 -8700 1078 -4900
rect 1238 -8700 1250 -4900
rect 1066 -8750 1250 -8700
rect 10750 -4900 10934 -4850
rect 10750 -8700 10762 -4900
rect 10922 -8700 10934 -4900
rect 10750 -8750 10934 -8700
rect 1066 -8762 10934 -8750
rect 1066 -8922 1300 -8762
rect 10700 -8922 10934 -8762
rect 1066 -8934 10934 -8922
<< mvpsubdiffcont >>
rect 1300 -238 10700 -78
rect 1078 -4100 1238 -300
rect 10762 -4100 10922 -300
rect 1300 -4322 10700 -4162
<< mvnsubdiffcont >>
rect 1300 -4838 10700 -4678
rect 1078 -8700 1238 -4900
rect 10762 -8700 10922 -4900
rect 1300 -8922 10700 -8762
<< locali >>
rect 1078 -300 1238 -78
rect -988 -4169 -760 -4135
rect 1078 -4322 1238 -4100
rect 10762 -300 10922 -78
rect 10762 -4322 10922 -4100
rect -2061 -4476 -2019 -4462
rect -2061 -4525 -2047 -4476
rect -1775 -4502 -1731 -4468
rect -1013 -4492 -896 -4462
rect -2061 -4539 -2019 -4525
rect -1013 -4542 -972 -4492
rect -922 -4542 -896 -4492
rect -1013 -4572 -896 -4542
rect 1078 -4900 1238 -4678
rect -988 -4983 -760 -4949
rect 1078 -8922 1238 -8700
rect 10762 -4900 10922 -4678
rect 10762 -8922 10922 -8700
<< viali >>
rect 1238 -238 1300 -78
rect 1300 -238 10700 -78
rect 10700 -238 10762 -78
rect 1078 -3966 1238 -434
rect -537 -4354 -503 -4320
rect 10762 -3966 10922 -434
rect 1238 -4322 1300 -4162
rect 1300 -4322 10700 -4162
rect 10700 -4322 10762 -4162
rect -2047 -4525 -1998 -4476
rect -2697 -4577 -2647 -4527
rect -2593 -4577 -2543 -4527
rect -2489 -4577 -2439 -4527
rect -972 -4542 -922 -4492
rect -249 -4502 -215 -4468
rect 1238 -4838 1300 -4678
rect 1300 -4838 10700 -4678
rect 10700 -4838 10762 -4678
rect 1078 -8566 1238 -5034
rect 10762 -8566 10922 -5034
rect 1238 -8922 1300 -8762
rect 1300 -8922 10700 -8762
rect 10700 -8922 10762 -8762
<< metal1 >>
rect -3087 141 -2313 147
rect -3087 -621 -3081 141
rect -2319 -621 -2313 141
rect -3087 -4129 -2313 -621
rect -1597 -19 -823 -13
rect -1597 -781 -1591 -19
rect -829 -781 -823 -19
rect -1597 -4129 -823 -781
rect -107 -19 667 -13
rect -107 -781 -101 -19
rect 661 -781 667 -19
rect -107 -4129 667 -781
rect 1072 -78 10928 -72
rect 1072 -238 1238 -78
rect 10762 -238 10928 -78
rect 1072 -244 10928 -238
rect 1072 -434 1244 -244
rect 1072 -3966 1078 -434
rect 1238 -738 1244 -434
rect 1844 -544 1854 -244
rect 10146 -544 10156 -244
rect 10756 -434 10928 -244
rect 10756 -738 10762 -434
rect 1238 -802 5765 -738
rect 1238 -2446 1244 -802
rect 4171 -1000 4217 -802
rect 4687 -1000 4733 -802
rect 5203 -1000 5249 -802
rect 5461 -836 5525 -830
rect 5461 -888 5467 -836
rect 5519 -888 5525 -836
rect 5461 -894 5525 -888
rect 5461 -1000 5507 -894
rect 5719 -1000 5765 -802
rect 6235 -802 10762 -738
rect 6235 -1000 6281 -802
rect 6475 -836 6539 -830
rect 6475 -888 6481 -836
rect 6533 -888 6539 -836
rect 6475 -894 6539 -888
rect 6493 -1000 6539 -894
rect 6751 -1000 6797 -802
rect 7267 -1000 7313 -802
rect 7783 -1000 7829 -802
rect 3655 -2032 3701 -2000
rect 3913 -2032 3959 -2000
rect 4429 -2032 4475 -2000
rect 4945 -2032 4991 -2000
rect 5977 -2032 6023 -2000
rect 7009 -2032 7055 -2000
rect 7525 -2032 7571 -2000
rect 8041 -2032 8087 -2000
rect 8299 -2032 8345 -2000
rect 3655 -2112 5143 -2032
rect 3655 -2164 3919 -2112
rect 3971 -2164 4025 -2112
rect 4105 -2164 4283 -2112
rect 4363 -2164 4426 -2112
rect 4478 -2164 4541 -2112
rect 4621 -2164 4799 -2112
rect 4879 -2164 4942 -2112
rect 4994 -2164 5057 -2112
rect 5137 -2164 5143 -2112
rect 3655 -2170 5143 -2164
rect 5309 -2112 5401 -2032
rect 5309 -2164 5315 -2112
rect 5395 -2164 5401 -2112
rect 5309 -2170 5401 -2164
rect 5567 -2112 5659 -2032
rect 5567 -2164 5573 -2112
rect 5653 -2164 5659 -2112
rect 5567 -2170 5659 -2164
rect 5825 -2112 6175 -2032
rect 5825 -2164 5831 -2112
rect 5911 -2126 6089 -2112
rect 5911 -2164 5969 -2126
rect 5825 -2170 5969 -2164
rect 1238 -2510 5507 -2446
rect 5963 -2488 5969 -2170
rect 6031 -2164 6089 -2126
rect 6169 -2164 6175 -2112
rect 6031 -2170 6175 -2164
rect 6341 -2112 6433 -2032
rect 6341 -2164 6347 -2112
rect 6427 -2164 6433 -2112
rect 6341 -2170 6433 -2164
rect 6599 -2112 6691 -2032
rect 6599 -2164 6605 -2112
rect 6685 -2164 6691 -2112
rect 6599 -2170 6691 -2164
rect 6857 -2112 8345 -2032
rect 6857 -2164 6863 -2112
rect 6943 -2164 7006 -2112
rect 7058 -2164 7121 -2112
rect 7201 -2164 7379 -2112
rect 7459 -2164 7522 -2112
rect 7574 -2164 7637 -2112
rect 7717 -2164 7895 -2112
rect 7975 -2164 8029 -2112
rect 8081 -2164 8345 -2112
rect 6857 -2170 8345 -2164
rect 6031 -2488 6037 -2170
rect 10756 -2446 10762 -802
rect 5963 -2494 6037 -2488
rect 1238 -3966 1244 -2510
rect 2365 -2722 2411 -2510
rect 2107 -2768 2213 -2722
rect 2305 -2768 2411 -2722
rect 2471 -2544 2563 -2538
rect 2471 -2596 2477 -2544
rect 2557 -2596 2563 -2544
rect 2471 -2768 2563 -2596
rect 3245 -2544 3337 -2538
rect 3245 -2596 3251 -2544
rect 3331 -2596 3337 -2544
rect 2623 -2636 2687 -2630
rect 2623 -2688 2629 -2636
rect 2681 -2688 2687 -2636
rect 2623 -2694 2687 -2688
rect 3130 -2636 3194 -2630
rect 3130 -2688 3136 -2636
rect 3188 -2688 3194 -2636
rect 3130 -2694 3194 -2688
rect 2107 -2800 2153 -2768
rect 2365 -2800 2411 -2768
rect 2623 -2800 2669 -2694
rect 3139 -2800 3185 -2694
rect 3245 -2768 3337 -2596
rect 3397 -2800 3443 -2510
rect 3503 -2544 3595 -2538
rect 3503 -2596 3509 -2544
rect 3589 -2596 3595 -2544
rect 3503 -2768 3595 -2596
rect 4277 -2544 4369 -2538
rect 4277 -2596 4283 -2544
rect 4363 -2596 4369 -2544
rect 3646 -2636 3710 -2630
rect 3646 -2688 3652 -2636
rect 3704 -2688 3710 -2636
rect 3646 -2694 3710 -2688
rect 4162 -2636 4226 -2630
rect 4162 -2688 4168 -2636
rect 4220 -2688 4226 -2636
rect 4162 -2694 4226 -2688
rect 3655 -2800 3701 -2694
rect 4171 -2800 4217 -2694
rect 4277 -2768 4369 -2596
rect 4429 -2800 4475 -2510
rect 4535 -2544 4627 -2538
rect 4535 -2596 4541 -2544
rect 4621 -2596 4627 -2544
rect 4535 -2768 4627 -2596
rect 5309 -2544 5401 -2538
rect 5309 -2596 5315 -2544
rect 5395 -2596 5401 -2544
rect 4678 -2636 4742 -2630
rect 4678 -2688 4684 -2636
rect 4736 -2688 4742 -2636
rect 4678 -2694 4742 -2688
rect 5194 -2636 5258 -2630
rect 5194 -2688 5200 -2636
rect 5252 -2688 5258 -2636
rect 5194 -2694 5258 -2688
rect 4687 -2800 4733 -2694
rect 5203 -2800 5249 -2694
rect 5309 -2768 5401 -2596
rect 5461 -2800 5507 -2510
rect 5567 -2544 5659 -2538
rect 5567 -2596 5573 -2544
rect 5653 -2596 5659 -2544
rect 5567 -2768 5659 -2596
rect 5968 -2544 6032 -2494
rect 6493 -2510 10762 -2446
rect 5968 -2596 5974 -2544
rect 6026 -2596 6032 -2544
rect 5968 -2602 6032 -2596
rect 6341 -2544 6433 -2538
rect 6341 -2596 6347 -2544
rect 6427 -2596 6433 -2544
rect 5710 -2636 5774 -2630
rect 5710 -2688 5716 -2636
rect 5768 -2688 5774 -2636
rect 5710 -2694 5774 -2688
rect 6226 -2636 6290 -2630
rect 6226 -2688 6232 -2636
rect 6284 -2688 6290 -2636
rect 6226 -2694 6290 -2688
rect 5719 -2800 5765 -2694
rect 6235 -2800 6281 -2694
rect 6341 -2768 6433 -2596
rect 6493 -2800 6539 -2510
rect 6599 -2544 6691 -2538
rect 6599 -2596 6605 -2544
rect 6685 -2596 6691 -2544
rect 6599 -2768 6691 -2596
rect 7373 -2544 7465 -2538
rect 7373 -2596 7379 -2544
rect 7459 -2596 7465 -2544
rect 6742 -2636 6806 -2630
rect 6742 -2688 6748 -2636
rect 6800 -2688 6806 -2636
rect 6742 -2694 6806 -2688
rect 7258 -2636 7322 -2630
rect 7258 -2688 7264 -2636
rect 7316 -2688 7322 -2636
rect 7258 -2694 7322 -2688
rect 6751 -2800 6797 -2694
rect 7267 -2800 7313 -2694
rect 7373 -2768 7465 -2596
rect 7525 -2800 7571 -2510
rect 7631 -2544 7723 -2538
rect 7631 -2596 7637 -2544
rect 7717 -2596 7723 -2544
rect 7631 -2768 7723 -2596
rect 8405 -2544 8497 -2538
rect 8405 -2596 8411 -2544
rect 8491 -2596 8497 -2544
rect 7774 -2636 7838 -2630
rect 7774 -2688 7780 -2636
rect 7832 -2688 7838 -2636
rect 7774 -2694 7838 -2688
rect 8290 -2636 8354 -2630
rect 8290 -2688 8296 -2636
rect 8348 -2688 8354 -2636
rect 8290 -2694 8354 -2688
rect 7783 -2800 7829 -2694
rect 8299 -2800 8345 -2694
rect 8405 -2768 8497 -2596
rect 8557 -2800 8603 -2510
rect 8663 -2544 8755 -2538
rect 8663 -2596 8669 -2544
rect 8749 -2596 8755 -2544
rect 8663 -2768 8755 -2596
rect 9437 -2544 9529 -2538
rect 9437 -2596 9443 -2544
rect 9523 -2596 9529 -2544
rect 8806 -2636 8870 -2630
rect 8806 -2688 8812 -2636
rect 8864 -2688 8870 -2636
rect 8806 -2694 8870 -2688
rect 9313 -2636 9377 -2630
rect 9313 -2688 9319 -2636
rect 9371 -2688 9377 -2636
rect 9313 -2694 9377 -2688
rect 8815 -2800 8861 -2694
rect 9331 -2800 9377 -2694
rect 9437 -2768 9529 -2596
rect 9589 -2722 9635 -2510
rect 9589 -2768 9695 -2722
rect 9787 -2768 9893 -2722
rect 9589 -2800 9635 -2768
rect 9847 -2800 9893 -2768
rect -3100 -4277 680 -4129
rect 1072 -4156 1244 -3966
rect 1844 -4156 1854 -3856
rect 2729 -4004 2821 -3878
rect 2881 -3906 2927 -3800
rect 2881 -3912 2945 -3906
rect 2881 -3964 2887 -3912
rect 2939 -3964 2945 -3912
rect 2881 -3970 2945 -3964
rect 2729 -4056 2735 -4004
rect 2815 -4056 2821 -4004
rect 2729 -4062 2821 -4056
rect 2987 -4004 3079 -3878
rect 2987 -4056 2993 -4004
rect 3073 -4056 3079 -4004
rect 2987 -4062 3079 -4056
rect 3761 -4004 3853 -3878
rect 3913 -3906 3959 -3800
rect 3904 -3912 3968 -3906
rect 3904 -3964 3910 -3912
rect 3962 -3964 3968 -3912
rect 3904 -3970 3968 -3964
rect 3761 -4056 3767 -4004
rect 3847 -4056 3853 -4004
rect 3761 -4062 3853 -4056
rect 4019 -4004 4111 -3878
rect 4019 -4056 4025 -4004
rect 4105 -4056 4111 -4004
rect 4019 -4062 4111 -4056
rect 4793 -4004 4885 -3878
rect 4945 -3906 4991 -3800
rect 4936 -3912 5000 -3906
rect 4936 -3964 4942 -3912
rect 4994 -3964 5000 -3912
rect 4936 -3970 5000 -3964
rect 4793 -4056 4799 -4004
rect 4879 -4056 4885 -4004
rect 4793 -4062 4885 -4056
rect 5051 -4004 5143 -3878
rect 5051 -4056 5057 -4004
rect 5137 -4056 5143 -4004
rect 5051 -4062 5143 -4056
rect 5825 -4004 5917 -3878
rect 5977 -3906 6023 -3800
rect 5968 -3912 6032 -3906
rect 5968 -3964 5974 -3912
rect 6026 -3964 6032 -3912
rect 5968 -3970 6032 -3964
rect 5825 -4056 5831 -4004
rect 5911 -4056 5917 -4004
rect 5825 -4062 5917 -4056
rect 5977 -4064 6023 -3970
rect 6083 -4004 6175 -3878
rect 6083 -4056 6089 -4004
rect 6169 -4056 6175 -4004
rect 6083 -4062 6175 -4056
rect 6857 -4004 6949 -3878
rect 7009 -3906 7055 -3800
rect 7000 -3912 7064 -3906
rect 7000 -3964 7006 -3912
rect 7058 -3964 7064 -3912
rect 7000 -3970 7064 -3964
rect 6857 -4056 6863 -4004
rect 6943 -4056 6949 -4004
rect 6857 -4062 6949 -4056
rect 7115 -4004 7207 -3878
rect 7115 -4056 7121 -4004
rect 7201 -4056 7207 -4004
rect 7115 -4062 7207 -4056
rect 7889 -4004 7981 -3878
rect 8041 -3906 8087 -3800
rect 8032 -3912 8096 -3906
rect 8032 -3964 8038 -3912
rect 8090 -3964 8096 -3912
rect 8032 -3970 8096 -3964
rect 7889 -4056 7895 -4004
rect 7975 -4056 7981 -4004
rect 7889 -4062 7981 -4056
rect 8147 -4004 8239 -3878
rect 8147 -4056 8153 -4004
rect 8233 -4056 8239 -4004
rect 8147 -4062 8239 -4056
rect 8921 -4004 9013 -3878
rect 9073 -3906 9119 -3800
rect 9055 -3912 9119 -3906
rect 9055 -3964 9061 -3912
rect 9113 -3964 9119 -3912
rect 9055 -3970 9119 -3964
rect 8921 -4056 8927 -4004
rect 9007 -4056 9013 -4004
rect 8921 -4062 9013 -4056
rect 9179 -4004 9271 -3878
rect 9179 -4056 9185 -4004
rect 9265 -4056 9271 -4004
rect 9179 -4062 9271 -4056
rect 5968 -4070 6032 -4064
rect 5968 -4122 5974 -4070
rect 6026 -4122 6032 -4070
rect 5968 -4128 6032 -4122
rect 10146 -4156 10156 -3856
rect 10756 -3966 10762 -2510
rect 10922 -3966 10928 -434
rect 10756 -4156 10928 -3966
rect 1072 -4162 10928 -4156
rect -549 -4320 -389 -4314
rect -549 -4354 -537 -4320
rect -503 -4354 -389 -4320
rect 1072 -4322 1238 -4162
rect 10762 -4322 10928 -4162
rect 1072 -4328 10928 -4322
rect -549 -4360 -389 -4354
rect -435 -4366 -389 -4360
rect -435 -4412 771 -4366
rect -2059 -4469 -1985 -4463
rect -2709 -4521 -2635 -4515
rect -2709 -4583 -2703 -4521
rect -2641 -4583 -2635 -4521
rect -2709 -4589 -2635 -4583
rect -2605 -4521 -2531 -4515
rect -2605 -4583 -2599 -4521
rect -2537 -4583 -2531 -4521
rect -2605 -4589 -2531 -4583
rect -2501 -4521 -2427 -4515
rect -2501 -4583 -2495 -4521
rect -2433 -4583 -2427 -4521
rect -2059 -4531 -2053 -4469
rect -1991 -4531 -1985 -4469
rect -753 -4468 -203 -4462
rect -2059 -4537 -1985 -4531
rect -984 -4486 -910 -4480
rect -984 -4548 -978 -4486
rect -916 -4496 -910 -4486
rect -753 -4496 -249 -4468
rect -916 -4502 -249 -4496
rect -215 -4502 -203 -4468
rect -916 -4508 -203 -4502
rect -916 -4542 -707 -4508
rect -916 -4548 -910 -4542
rect -984 -4554 -910 -4548
rect -2501 -4589 -2427 -4583
rect 725 -4565 771 -4412
rect 875 -4565 881 -4562
rect 725 -4611 881 -4565
rect 875 -4614 881 -4611
rect 933 -4614 939 -4562
rect 1072 -4678 10928 -4672
rect 1072 -4838 1238 -4678
rect 10762 -4838 10928 -4678
rect -3100 -4989 680 -4841
rect 1072 -4844 10928 -4838
rect -3087 -8219 -2313 -4989
rect -3087 -8981 -3081 -8219
rect -2319 -8981 -2313 -8219
rect -3087 -8987 -2313 -8981
rect -1597 -8219 -823 -4989
rect -1597 -8981 -1591 -8219
rect -829 -8981 -823 -8219
rect -1597 -8987 -823 -8981
rect -107 -8219 667 -4989
rect -107 -8981 -101 -8219
rect 661 -8981 667 -8219
rect 1072 -5034 1244 -4844
rect 1072 -8566 1078 -5034
rect 1238 -6730 1244 -5034
rect 1844 -5144 1854 -4844
rect 5968 -4878 6032 -4872
rect 5968 -4930 5974 -4878
rect 6026 -4930 6032 -4878
rect 5968 -4936 6032 -4930
rect 5825 -5027 5917 -5021
rect 5825 -5079 5831 -5027
rect 5911 -5079 5917 -5027
rect 5825 -5159 5917 -5079
rect 5977 -5200 6023 -4936
rect 6083 -5027 6175 -5021
rect 6083 -5079 6089 -5027
rect 6169 -5079 6175 -5027
rect 6083 -5159 6175 -5079
rect 10146 -5144 10156 -4844
rect 10756 -5034 10928 -4844
rect 5461 -6241 5507 -6200
rect 5719 -6241 5765 -6200
rect 5461 -6287 5765 -6241
rect 5719 -6306 5765 -6287
rect 6235 -6241 6281 -6200
rect 6493 -6241 6539 -6200
rect 6235 -6287 6539 -6241
rect 6235 -6306 6281 -6287
rect 5719 -6312 5783 -6306
rect 5719 -6364 5725 -6312
rect 5777 -6364 5783 -6312
rect 5719 -6370 5783 -6364
rect 5968 -6312 6032 -6306
rect 5968 -6364 5974 -6312
rect 6026 -6364 6032 -6312
rect 1238 -6794 5894 -6730
rect 1238 -8566 1244 -6794
rect 4816 -6913 4862 -6794
rect 4558 -7000 4862 -6913
rect 5332 -7000 5378 -6794
rect 5590 -6836 5654 -6830
rect 5590 -6888 5596 -6836
rect 5648 -6888 5654 -6836
rect 5590 -6894 5654 -6888
rect 5590 -7000 5636 -6894
rect 5848 -6913 5894 -6794
rect 5968 -6827 6032 -6364
rect 6217 -6312 6281 -6306
rect 6217 -6364 6223 -6312
rect 6275 -6364 6281 -6312
rect 6217 -6370 6281 -6364
rect 10756 -6730 10762 -5034
rect 5968 -6879 5974 -6827
rect 6026 -6879 6032 -6827
rect 6622 -6794 10762 -6730
rect 5968 -6885 6032 -6879
rect 6346 -6836 6410 -6830
rect 6346 -6888 6352 -6836
rect 6404 -6888 6410 -6836
rect 6346 -6894 6410 -6888
rect 5696 -7000 5894 -6913
rect 6212 -6922 6318 -6913
rect 6364 -6922 6410 -6894
rect 6212 -7000 6410 -6922
rect 6622 -7000 6668 -6794
rect 7138 -6913 7184 -6794
rect 7138 -7000 7442 -6913
rect 5074 -8041 5120 -8000
rect 6106 -8041 6152 -8000
rect 6880 -8041 6926 -8000
rect 4922 -8112 5272 -8041
rect 4922 -8164 4928 -8112
rect 5008 -8164 5071 -8112
rect 5123 -8164 5186 -8112
rect 5266 -8164 5272 -8112
rect 4922 -8170 5272 -8164
rect 5438 -8112 5530 -8041
rect 5438 -8164 5444 -8112
rect 5524 -8164 5530 -8112
rect 5438 -8170 5530 -8164
rect 5954 -8112 6161 -8041
rect 5954 -8164 5960 -8112
rect 6040 -8164 6103 -8112
rect 6155 -8164 6161 -8112
rect 5954 -8170 6161 -8164
rect 6470 -8112 6562 -8041
rect 6470 -8164 6476 -8112
rect 6556 -8164 6562 -8112
rect 6470 -8170 6562 -8164
rect 6728 -8112 7078 -8041
rect 6728 -8164 6734 -8112
rect 6814 -8164 6877 -8112
rect 6929 -8164 6992 -8112
rect 7072 -8164 7078 -8112
rect 6728 -8170 7078 -8164
rect 1072 -8756 1244 -8566
rect 1844 -8756 1854 -8456
rect 10146 -8756 10156 -8456
rect 10756 -8566 10762 -6794
rect 10922 -8566 10928 -5034
rect 10756 -8756 10928 -8566
rect 1072 -8762 10928 -8756
rect 1072 -8922 1238 -8762
rect 10762 -8922 10928 -8762
rect 1072 -8928 10928 -8922
rect -107 -8987 667 -8981
<< via1 >>
rect -3081 -621 -2319 141
rect -1591 -781 -829 -19
rect -101 -781 661 -19
rect 1244 -544 1844 -244
rect 10156 -544 10756 -244
rect 5467 -888 5519 -836
rect 6481 -888 6533 -836
rect 3919 -2164 3971 -2112
rect 4025 -2164 4105 -2112
rect 4283 -2164 4363 -2112
rect 4426 -2164 4478 -2112
rect 4541 -2164 4621 -2112
rect 4799 -2164 4879 -2112
rect 4942 -2164 4994 -2112
rect 5057 -2164 5137 -2112
rect 5315 -2164 5395 -2112
rect 5573 -2164 5653 -2112
rect 5831 -2164 5911 -2112
rect 5969 -2488 6031 -2126
rect 6089 -2164 6169 -2112
rect 6347 -2164 6427 -2112
rect 6605 -2164 6685 -2112
rect 6863 -2164 6943 -2112
rect 7006 -2164 7058 -2112
rect 7121 -2164 7201 -2112
rect 7379 -2164 7459 -2112
rect 7522 -2164 7574 -2112
rect 7637 -2164 7717 -2112
rect 7895 -2164 7975 -2112
rect 8029 -2164 8081 -2112
rect 2477 -2596 2557 -2544
rect 3251 -2596 3331 -2544
rect 2629 -2688 2681 -2636
rect 3136 -2688 3188 -2636
rect 3509 -2596 3589 -2544
rect 4283 -2596 4363 -2544
rect 3652 -2688 3704 -2636
rect 4168 -2688 4220 -2636
rect 4541 -2596 4621 -2544
rect 5315 -2596 5395 -2544
rect 4684 -2688 4736 -2636
rect 5200 -2688 5252 -2636
rect 5573 -2596 5653 -2544
rect 5974 -2596 6026 -2544
rect 6347 -2596 6427 -2544
rect 5716 -2688 5768 -2636
rect 6232 -2688 6284 -2636
rect 6605 -2596 6685 -2544
rect 7379 -2596 7459 -2544
rect 6748 -2688 6800 -2636
rect 7264 -2688 7316 -2636
rect 7637 -2596 7717 -2544
rect 8411 -2596 8491 -2544
rect 7780 -2688 7832 -2636
rect 8296 -2688 8348 -2636
rect 8669 -2596 8749 -2544
rect 9443 -2596 9523 -2544
rect 8812 -2688 8864 -2636
rect 9319 -2688 9371 -2636
rect 1244 -4156 1844 -3856
rect 2887 -3964 2939 -3912
rect 2735 -4056 2815 -4004
rect 2993 -4056 3073 -4004
rect 3910 -3964 3962 -3912
rect 3767 -4056 3847 -4004
rect 4025 -4056 4105 -4004
rect 4942 -3964 4994 -3912
rect 4799 -4056 4879 -4004
rect 5057 -4056 5137 -4004
rect 5974 -3964 6026 -3912
rect 5831 -4056 5911 -4004
rect 6089 -4056 6169 -4004
rect 7006 -3964 7058 -3912
rect 6863 -4056 6943 -4004
rect 7121 -4056 7201 -4004
rect 8038 -3964 8090 -3912
rect 7895 -4056 7975 -4004
rect 8153 -4056 8233 -4004
rect 9061 -3964 9113 -3912
rect 8927 -4056 9007 -4004
rect 9185 -4056 9265 -4004
rect 5974 -4122 6026 -4070
rect 10156 -4156 10756 -3856
rect -2703 -4527 -2641 -4521
rect -2703 -4577 -2697 -4527
rect -2697 -4577 -2647 -4527
rect -2647 -4577 -2641 -4527
rect -2703 -4583 -2641 -4577
rect -2599 -4527 -2537 -4521
rect -2599 -4577 -2593 -4527
rect -2593 -4577 -2543 -4527
rect -2543 -4577 -2537 -4527
rect -2599 -4583 -2537 -4577
rect -2495 -4527 -2433 -4521
rect -2495 -4577 -2489 -4527
rect -2489 -4577 -2439 -4527
rect -2439 -4577 -2433 -4527
rect -2495 -4583 -2433 -4577
rect -2053 -4476 -1991 -4469
rect -2053 -4525 -2047 -4476
rect -2047 -4525 -1998 -4476
rect -1998 -4525 -1991 -4476
rect -2053 -4531 -1991 -4525
rect -978 -4492 -916 -4486
rect -978 -4542 -972 -4492
rect -972 -4542 -922 -4492
rect -922 -4542 -916 -4492
rect -978 -4548 -916 -4542
rect 881 -4614 933 -4562
rect -3081 -8981 -2319 -8219
rect -1591 -8981 -829 -8219
rect -101 -8981 661 -8219
rect 1244 -5144 1844 -4844
rect 5974 -4930 6026 -4878
rect 5831 -5079 5911 -5027
rect 6089 -5079 6169 -5027
rect 10156 -5144 10756 -4844
rect 5725 -6364 5777 -6312
rect 5974 -6364 6026 -6312
rect 5596 -6888 5648 -6836
rect 6223 -6364 6275 -6312
rect 5974 -6879 6026 -6827
rect 6352 -6888 6404 -6836
rect 4928 -8164 5008 -8112
rect 5071 -8164 5123 -8112
rect 5186 -8164 5266 -8112
rect 5444 -8164 5524 -8112
rect 5960 -8164 6040 -8112
rect 6103 -8164 6155 -8112
rect 6476 -8164 6556 -8112
rect 6734 -8164 6814 -8112
rect 6877 -8164 6929 -8112
rect 6992 -8164 7072 -8112
rect 1244 -8756 1844 -8456
rect 10156 -8756 10756 -8456
<< metal2 >>
rect -3087 141 -2313 147
rect -3087 -621 -3081 141
rect -2319 -621 -2313 141
rect -3087 -627 -2313 -621
rect -1597 -19 -823 -13
rect -1597 -781 -1591 -19
rect -829 -781 -823 -19
rect -1597 -787 -823 -781
rect -107 -19 667 -13
rect -107 -781 -101 -19
rect 661 -781 667 -19
rect 1244 -244 1844 -230
rect 1244 -553 1844 -544
rect 10156 -244 10756 -230
rect 10156 -553 10756 -544
rect -107 -787 667 -781
rect 5968 -710 9991 -646
rect 5968 -830 6032 -710
rect 5461 -836 6539 -830
rect 5461 -888 5467 -836
rect 5519 -888 6481 -836
rect 6533 -888 6539 -836
rect 5461 -894 6539 -888
rect 3913 -2112 8087 -2106
rect 3913 -2164 3919 -2112
rect 3971 -2164 4025 -2112
rect 4105 -2164 4283 -2112
rect 4363 -2164 4426 -2112
rect 4478 -2164 4541 -2112
rect 4621 -2164 4799 -2112
rect 4879 -2164 4942 -2112
rect 4994 -2164 5057 -2112
rect 5137 -2164 5315 -2112
rect 5395 -2164 5573 -2112
rect 5653 -2164 5831 -2112
rect 5911 -2126 6089 -2112
rect 5911 -2164 5969 -2126
rect 3913 -2170 5969 -2164
rect 5963 -2488 5969 -2170
rect 6031 -2164 6089 -2126
rect 6169 -2164 6347 -2112
rect 6427 -2164 6605 -2112
rect 6685 -2164 6863 -2112
rect 6943 -2164 7006 -2112
rect 7058 -2164 7121 -2112
rect 7201 -2164 7379 -2112
rect 7459 -2164 7522 -2112
rect 7574 -2164 7637 -2112
rect 7717 -2164 7895 -2112
rect 7975 -2164 8029 -2112
rect 8081 -2164 8087 -2112
rect 6031 -2170 8087 -2164
rect 6031 -2488 6037 -2170
rect 5963 -2494 6037 -2488
rect 2471 -2544 9529 -2538
rect 2471 -2596 2477 -2544
rect 2557 -2596 3251 -2544
rect 3331 -2596 3509 -2544
rect 3589 -2596 4283 -2544
rect 4363 -2596 4541 -2544
rect 4621 -2596 5315 -2544
rect 5395 -2596 5573 -2544
rect 5653 -2596 5974 -2544
rect 6026 -2596 6347 -2544
rect 6427 -2596 6605 -2544
rect 6685 -2596 7379 -2544
rect 7459 -2596 7637 -2544
rect 7717 -2596 8411 -2544
rect 8491 -2596 8669 -2544
rect 8749 -2596 9443 -2544
rect 9523 -2596 9529 -2544
rect 2471 -2602 9529 -2596
rect 2623 -2636 9377 -2630
rect 2623 -2688 2629 -2636
rect 2681 -2688 3136 -2636
rect 3188 -2688 3652 -2636
rect 3704 -2688 4168 -2636
rect 4220 -2688 4684 -2636
rect 4736 -2688 5200 -2636
rect 5252 -2688 5716 -2636
rect 5768 -2688 6232 -2636
rect 6284 -2688 6748 -2636
rect 6800 -2688 7264 -2636
rect 7316 -2688 7780 -2636
rect 7832 -2688 8296 -2636
rect 8348 -2688 8812 -2636
rect 8864 -2688 9319 -2636
rect 9371 -2688 9377 -2636
rect 2623 -2694 9377 -2688
rect 1244 -3856 1844 -3846
rect 2881 -3912 9119 -3906
rect 2881 -3964 2887 -3912
rect 2939 -3964 3910 -3912
rect 3962 -3964 4942 -3912
rect 4994 -3964 5974 -3912
rect 6026 -3964 7006 -3912
rect 7058 -3964 8038 -3912
rect 8090 -3964 9061 -3912
rect 9113 -3964 9119 -3912
rect 2881 -3970 9119 -3964
rect 2729 -4004 9271 -3998
rect 2729 -4056 2735 -4004
rect 2815 -4056 2993 -4004
rect 3073 -4056 3767 -4004
rect 3847 -4056 4025 -4004
rect 4105 -4056 4799 -4004
rect 4879 -4056 5057 -4004
rect 5137 -4056 5831 -4004
rect 5911 -4031 6089 -4004
rect 5911 -4056 5935 -4031
rect 2729 -4062 5935 -4056
rect 6065 -4056 6089 -4031
rect 6169 -4056 6863 -4004
rect 6943 -4056 7121 -4004
rect 7201 -4056 7895 -4004
rect 7975 -4056 8153 -4004
rect 8233 -4056 8927 -4004
rect 9007 -4056 9185 -4004
rect 9265 -4056 9271 -4004
rect 1244 -4166 1844 -4156
rect -2059 -4469 -1985 -4463
rect -2709 -4521 -2635 -4515
rect -2709 -4583 -2703 -4521
rect -2641 -4583 -2635 -4521
rect -2709 -4589 -2635 -4583
rect -2605 -4521 -2531 -4515
rect -2605 -4583 -2599 -4521
rect -2537 -4583 -2531 -4521
rect -2605 -4589 -2531 -4583
rect -2501 -4521 -2427 -4515
rect -2501 -4583 -2495 -4521
rect -2433 -4583 -2427 -4521
rect -2059 -4531 -2053 -4469
rect -1991 -4531 -1985 -4469
rect -2059 -4537 -1985 -4531
rect -984 -4486 -910 -4480
rect -984 -4548 -978 -4486
rect -916 -4548 -910 -4486
rect 4420 -4506 4484 -4062
rect 5963 -4068 6037 -4059
rect 6065 -4062 9271 -4056
rect 5963 -4124 5972 -4068
rect 6028 -4124 6037 -4068
rect 5963 -4133 6037 -4124
rect 4415 -4515 4489 -4506
rect -984 -4554 -910 -4548
rect -2501 -4589 -2427 -4583
rect 848 -4624 866 -4524
rect 966 -4624 975 -4524
rect 4415 -4571 4424 -4515
rect 4480 -4571 4489 -4515
rect 4415 -4580 4489 -4571
rect 1244 -4844 1844 -4834
rect 4420 -5021 4484 -4580
rect 5968 -4878 6032 -4133
rect 7516 -4506 7580 -4062
rect 7511 -4515 7585 -4506
rect 7511 -4571 7520 -4515
rect 7576 -4571 7585 -4515
rect 7511 -4580 7585 -4571
rect 5968 -4930 5974 -4878
rect 6026 -4930 6032 -4878
rect 5968 -4936 6032 -4930
rect 7516 -5021 7580 -4580
rect 4420 -5027 7580 -5021
rect 4420 -5079 5831 -5027
rect 5911 -5079 6089 -5027
rect 6169 -5079 7580 -5027
rect 1244 -5154 1844 -5144
rect 5719 -6312 6281 -6306
rect 5719 -6364 5725 -6312
rect 5777 -6364 5974 -6312
rect 6026 -6364 6223 -6312
rect 6275 -6364 6281 -6312
rect 5719 -6370 6281 -6364
rect 5968 -6827 6032 -6822
rect 5968 -6830 5974 -6827
rect 5590 -6836 5974 -6830
rect 5590 -6888 5596 -6836
rect 5648 -6879 5974 -6836
rect 6026 -6830 6032 -6827
rect 6026 -6836 6410 -6830
rect 6026 -6879 6352 -6836
rect 5648 -6888 6352 -6879
rect 6404 -6888 6410 -6836
rect 5590 -6894 6410 -6888
rect 4922 -8112 7078 -8106
rect 4922 -8164 4928 -8112
rect 5008 -8164 5071 -8112
rect 5123 -8164 5186 -8112
rect 5266 -8164 5444 -8112
rect 5524 -8164 5960 -8112
rect 6040 -8164 6103 -8112
rect 6155 -8164 6476 -8112
rect 6556 -8164 6734 -8112
rect 6814 -8164 6877 -8112
rect 6929 -8164 6992 -8112
rect 7072 -8164 7078 -8112
rect 4922 -8170 7078 -8164
rect 5954 -8198 6046 -8170
rect 9927 -8198 9991 -710
rect 10156 -3856 10756 -3846
rect 10156 -4166 10756 -4156
rect 10156 -4844 10756 -4834
rect 10156 -5154 10756 -5144
rect -3087 -8219 -2313 -8213
rect -3087 -8981 -3081 -8219
rect -2319 -8981 -2313 -8219
rect -3087 -8987 -2313 -8981
rect -1597 -8219 -823 -8213
rect -1597 -8981 -1591 -8219
rect -829 -8981 -823 -8219
rect -1597 -8987 -823 -8981
rect -107 -8219 667 -8213
rect -107 -8981 -101 -8219
rect 661 -8981 667 -8219
rect 5954 -8262 9991 -8198
rect 1244 -8456 1844 -8442
rect 1244 -8765 1844 -8756
rect 10156 -8456 10756 -8442
rect 10156 -8765 10756 -8756
rect -107 -8987 667 -8981
<< via2 >>
rect -3078 -618 -2322 138
rect -1588 -778 -832 -22
rect -98 -778 658 -22
rect 1244 -544 1844 -244
rect 10156 -544 10756 -244
rect 5972 -2485 6028 -2129
rect 1244 -4156 1844 -3856
rect -2700 -4580 -2644 -4524
rect -2596 -4580 -2540 -4524
rect -2492 -4580 -2436 -4524
rect -2050 -4528 -1994 -4472
rect -975 -4545 -919 -4489
rect 5972 -4070 6028 -4068
rect 5972 -4122 5974 -4070
rect 5974 -4122 6026 -4070
rect 6026 -4122 6028 -4070
rect 5972 -4124 6028 -4122
rect 866 -4562 966 -4524
rect 866 -4614 881 -4562
rect 881 -4614 933 -4562
rect 933 -4614 966 -4562
rect 866 -4624 966 -4614
rect 4424 -4571 4480 -4515
rect 1244 -5144 1844 -4844
rect 7520 -4571 7576 -4515
rect 10156 -4156 10756 -3856
rect 10156 -5144 10756 -4844
rect -3078 -8978 -2322 -8222
rect -1588 -8978 -832 -8222
rect -98 -8978 658 -8222
rect 1244 -8756 1844 -8456
rect 10156 -8756 10756 -8456
<< metal3 >>
rect -10100 5900 -3500 8000
rect -3100 5900 3500 8000
rect 3900 7200 10500 8000
rect 10580 7900 11020 8000
rect 10580 7200 10680 7900
rect 3900 5900 10680 7200
rect -10740 5676 -10420 5736
rect -10740 3274 -10679 5676
rect -10479 5275 -10420 5676
rect -10100 5600 10680 5900
rect -10100 5275 10500 5600
rect -10479 4300 10500 5275
rect -10479 3675 -3500 4300
rect -10479 3274 -10420 3675
rect -10740 3214 -10420 3274
rect -10100 1800 -3500 3675
rect -3100 1800 3500 4300
rect 3900 4200 10500 4300
rect 10580 4200 10680 5600
rect 3900 2600 10680 4200
rect 3900 1800 10500 2600
rect 10580 1500 10680 2600
rect 10920 1500 11020 7900
rect 10580 1400 11020 1500
rect -3100 154 -2300 160
rect -3100 -634 -3094 154
rect -2306 -634 -2300 154
rect -3100 -640 -2300 -634
rect -1610 -6 -810 0
rect -10900 -1120 -2628 -720
rect -1610 -794 -1604 -6
rect -816 -794 -810 -6
rect -1610 -800 -810 -794
rect -120 -6 680 0
rect -120 -794 -114 -6
rect 674 -794 680 -6
rect 1234 -244 1854 -239
rect 1234 -544 1244 -244
rect 1844 -544 1854 -244
rect 1234 -549 1854 -544
rect 10146 -244 10766 -239
rect 10146 -544 10156 -244
rect 10756 -544 10766 -244
rect 10146 -549 10766 -544
rect -120 -800 680 -794
rect -10900 -4600 -10500 -1120
rect -12000 -5000 -10500 -4600
rect -10740 -5338 -10420 -5278
rect -10740 -7740 -10680 -5338
rect -10480 -5739 -10420 -5338
rect -10100 -5739 -3500 -1200
rect -3000 -2135 -2628 -1120
rect 5600 -2129 6050 -2107
rect 5600 -2135 5972 -2129
rect -3000 -2485 5972 -2135
rect 6028 -2485 6050 -2129
rect -3000 -2507 6050 -2485
rect -1410 -3431 -1010 -3371
rect -1410 -3671 -1350 -3431
rect -3284 -3711 -1350 -3671
rect -1070 -3671 -1010 -3431
rect -1070 -3711 2034 -3671
rect -3284 -3771 2034 -3711
rect -3284 -4502 -3184 -3771
rect 1234 -3856 1854 -3851
rect -997 -4096 965 -3996
rect -2072 -4472 -1972 -4450
rect -3284 -4524 -2414 -4502
rect -3284 -4580 -2700 -4524
rect -2644 -4580 -2596 -4524
rect -2540 -4580 -2492 -4524
rect -2436 -4580 -2414 -4524
rect -3284 -4602 -2414 -4580
rect -2072 -4528 -2050 -4472
rect -1994 -4528 -1972 -4472
rect -10480 -7339 -3500 -5739
rect -2072 -6400 -1972 -4528
rect -997 -4489 -897 -4096
rect 865 -4333 965 -4096
rect 1234 -4156 1244 -3856
rect 1844 -4156 1854 -3856
rect 1934 -4046 2034 -3771
rect 10146 -3856 10766 -3851
rect 1934 -4068 6050 -4046
rect 1934 -4124 5972 -4068
rect 6028 -4124 6050 -4068
rect 1934 -4146 6050 -4124
rect 1234 -4161 1854 -4156
rect 10146 -4156 10156 -3856
rect 10756 -4156 10766 -3856
rect 10146 -4161 10766 -4156
rect 10972 -4108 11983 -4008
rect 865 -4433 6050 -4333
rect 10972 -4405 11072 -4108
rect -997 -4545 -975 -4489
rect -919 -4545 -897 -4489
rect 5950 -4493 6050 -4433
rect 4402 -4515 7598 -4493
rect -997 -4567 -897 -4545
rect 861 -4524 971 -4519
rect 861 -4624 866 -4524
rect 966 -4624 4088 -4524
rect 4402 -4571 4424 -4515
rect 4480 -4571 7520 -4515
rect 7576 -4571 7598 -4515
rect 4402 -4593 7598 -4571
rect 9071 -4505 11072 -4405
rect 861 -4629 971 -4624
rect 3988 -4789 4088 -4624
rect 9071 -4789 9171 -4505
rect 1234 -4844 1854 -4839
rect 1234 -5144 1244 -4844
rect 1844 -5144 1854 -4844
rect 3988 -4889 9171 -4789
rect 10146 -4844 10766 -4839
rect 1234 -5149 1854 -5144
rect 10146 -5144 10156 -4844
rect 10756 -5144 10766 -4844
rect 10146 -5149 10766 -5144
rect 11200 -5000 12000 -4600
rect 11200 -6400 11600 -5000
rect -2072 -6800 11600 -6400
rect -10480 -7740 -10420 -7339
rect -10100 -7400 -3500 -7339
rect -10740 -7800 -10420 -7740
rect -3100 -8206 -2300 -8200
rect -3100 -8994 -3094 -8206
rect -2306 -8994 -2300 -8206
rect -3100 -9000 -2300 -8994
rect -1610 -8206 -810 -8200
rect -1610 -8994 -1604 -8206
rect -816 -8994 -810 -8206
rect -1610 -9000 -810 -8994
rect -120 -8206 680 -8200
rect -120 -8994 -114 -8206
rect 674 -8994 680 -8206
rect 1234 -8456 1854 -8451
rect 1234 -8756 1244 -8456
rect 1844 -8756 1854 -8456
rect 1234 -8761 1854 -8756
rect 10146 -8456 10766 -8451
rect 10146 -8756 10156 -8456
rect 10756 -8756 10766 -8456
rect 10146 -8761 10766 -8756
rect -120 -9000 680 -8994
<< via3 >>
rect -10679 3274 -10479 5676
rect 10680 1500 10920 7900
rect -3094 138 -2306 154
rect -3094 -618 -3078 138
rect -3078 -618 -2322 138
rect -2322 -618 -2306 138
rect -3094 -634 -2306 -618
rect -1604 -22 -816 -6
rect -1604 -778 -1588 -22
rect -1588 -778 -832 -22
rect -832 -778 -816 -22
rect -1604 -794 -816 -778
rect -114 -22 674 -6
rect -114 -778 -98 -22
rect -98 -778 658 -22
rect 658 -778 674 -22
rect -114 -794 674 -778
rect 1244 -544 1844 -244
rect 10156 -544 10756 -244
rect -10680 -7740 -10480 -5338
rect -1350 -3711 -1070 -3431
rect 1244 -4156 1844 -3856
rect 10156 -4156 10756 -3856
rect 1244 -5144 1844 -4844
rect 10156 -5144 10756 -4844
rect -3094 -8222 -2306 -8206
rect -3094 -8978 -3078 -8222
rect -3078 -8978 -2322 -8222
rect -2322 -8978 -2306 -8222
rect -3094 -8994 -2306 -8978
rect -1604 -8222 -816 -8206
rect -1604 -8978 -1588 -8222
rect -1588 -8978 -832 -8222
rect -832 -8978 -816 -8222
rect -1604 -8994 -816 -8978
rect -114 -8222 674 -8206
rect -114 -8978 -98 -8222
rect -98 -8978 658 -8222
rect 658 -8978 674 -8222
rect -114 -8994 674 -8978
rect 1244 -8756 1844 -8456
rect 10156 -8756 10756 -8456
<< mimcap >>
rect -10000 7850 -3600 7900
rect -10000 1950 -3950 7850
rect -3650 1950 -3600 7850
rect -10000 1900 -3600 1950
rect -3000 7850 3400 7900
rect -3000 1950 3050 7850
rect 3350 1950 3400 7850
rect -3000 1900 3400 1950
rect 4000 7850 10400 7900
rect 4000 1950 10050 7850
rect 10350 1950 10400 7850
rect 4000 1900 10400 1950
rect -10000 -1350 -3600 -1300
rect -10000 -7250 -3950 -1350
rect -3650 -7250 -3600 -1350
rect -10000 -7300 -3600 -7250
<< mimcapcontact >>
rect -3950 1950 -3650 7850
rect 3050 1950 3350 7850
rect 10050 1950 10350 7850
rect -3950 -7250 -3650 -1350
<< metal4 >>
rect -12000 8900 12000 9000
rect -12000 8300 -11800 8900
rect -11200 8300 12000 8900
rect -12000 8200 12000 8300
rect -10100 7850 -3500 8000
rect -10740 5676 -10420 5736
rect -10740 3274 -10697 5676
rect -10461 3274 -10420 5676
rect -10740 3214 -10420 3274
rect -10100 1950 -3950 7850
rect -3650 1950 -3500 7850
rect -10100 1800 -3500 1950
rect -3100 7850 3500 8000
rect -3100 1950 3050 7850
rect 3350 1950 3500 7850
rect -3100 1800 3500 1950
rect 3900 7850 10500 8000
rect 3900 1950 10050 7850
rect 10350 1950 10500 7850
rect 3900 1800 10500 1950
rect 10580 7900 11020 8000
rect -10100 1400 -3900 1800
rect -3100 1400 3100 1800
rect 3900 1400 10100 1800
rect 10580 1500 10680 7900
rect 10920 1500 11020 7900
rect 10580 1400 11020 1500
rect -7700 800 -6100 1400
rect -700 800 900 1400
rect 6300 800 7900 1400
rect -12000 154 12000 800
rect -12000 -634 -3094 154
rect -2306 -6 12000 154
rect -2306 -634 -1604 -6
rect -12000 -794 -1604 -634
rect -816 -794 -114 -6
rect 674 -244 12000 -6
rect 674 -544 1244 -244
rect 1844 -544 10156 -244
rect 10756 -544 12000 -244
rect 674 -794 12000 -544
rect -12000 -800 12000 -794
rect -7700 -1200 -6100 -800
rect -10100 -1350 -3500 -1200
rect -10740 -5338 -10420 -5278
rect -10740 -7740 -10698 -5338
rect -10462 -7740 -10420 -5338
rect -10740 -7800 -10420 -7740
rect -10100 -7250 -3950 -1350
rect -3650 -7250 -3500 -1350
rect -1410 -3431 -1010 -3371
rect -1410 -3711 -1350 -3431
rect -1070 -3711 -1010 -3431
rect -1410 -3771 -1010 -3711
rect 1243 -3856 1845 -3855
rect 1243 -4156 1244 -3856
rect 1844 -4156 1845 -3856
rect 1243 -4157 1845 -4156
rect 10155 -3856 10757 -3855
rect 10155 -4156 10156 -3856
rect 10756 -4156 10757 -3856
rect 10155 -4157 10757 -4156
rect 1243 -4844 1845 -4843
rect 1243 -5144 1244 -4844
rect 1844 -5144 1845 -4844
rect 1243 -5145 1845 -5144
rect 10155 -4844 10757 -4843
rect 10155 -5144 10156 -4844
rect 10756 -5144 10757 -4844
rect 10155 -5145 10757 -5144
rect -10100 -7400 -3500 -7250
rect -10100 -7800 -3900 -7400
rect -12000 -8206 12000 -8200
rect -12000 -8300 -3094 -8206
rect -12000 -8900 -11800 -8300
rect -11200 -8900 -3094 -8300
rect -12000 -8994 -3094 -8900
rect -2306 -8994 -1604 -8206
rect -816 -8994 -114 -8206
rect 674 -8456 12000 -8206
rect 674 -8756 1244 -8456
rect 1844 -8756 10156 -8456
rect 10756 -8756 12000 -8456
rect 674 -8994 12000 -8756
rect -12000 -9000 12000 -8994
<< via4 >>
rect -11800 8300 -11200 8900
rect -10697 3274 -10679 5676
rect -10679 3274 -10479 5676
rect -10479 3274 -10461 5676
rect 10680 1500 10920 7900
rect -10698 -7740 -10680 -5338
rect -10680 -7740 -10480 -5338
rect -10480 -7740 -10462 -5338
rect -1350 -3711 -1070 -3431
rect -11800 -8900 -11200 -8300
<< mimcap2 >>
rect -10000 1850 -4000 7900
rect -10000 1550 -9950 1850
rect -4050 1550 -4000 1850
rect -10000 1500 -4000 1550
rect -3000 1850 3000 7900
rect -3000 1550 -2950 1850
rect 2950 1550 3000 1850
rect -3000 1500 3000 1550
rect 4000 1850 10000 7900
rect 4000 1550 4050 1850
rect 9950 1550 10000 1850
rect 4000 1500 10000 1550
rect -10000 -7350 -4000 -1300
rect -10000 -7650 -9950 -7350
rect -4050 -7650 -4000 -7350
rect -10000 -7700 -4000 -7650
<< mimcap2contact >>
rect -9950 1550 -4050 1850
rect -2950 1550 2950 1850
rect 4050 1550 9950 1850
rect -9950 -7650 -4050 -7350
<< metal5 >>
rect -12000 8900 -11000 9000
rect -12000 8300 -11800 8900
rect -11200 8300 -11000 8900
rect -12000 6056 -11000 8300
rect -12000 2894 -11060 6056
rect -10100 5900 -3900 8000
rect -3100 5900 3100 8000
rect 3900 6800 10100 8000
rect 10580 7900 11020 8000
rect 10580 6800 10680 7900
rect 3900 5900 10680 6800
rect -10740 5676 -10420 5736
rect -10740 3274 -10697 5676
rect -10461 5275 -10420 5676
rect -10100 5275 10680 5900
rect -10461 5200 10680 5275
rect -10461 4300 10100 5200
rect -10461 3675 -3900 4300
rect -10461 3274 -10420 3675
rect -10740 3214 -10420 3274
rect -12000 -4958 -11000 2894
rect -10100 1850 -3900 3675
rect -10100 1550 -9950 1850
rect -4050 1550 -3900 1850
rect -10100 1400 -3900 1550
rect -3100 1850 3100 4300
rect -3100 1550 -2950 1850
rect 2950 1550 3100 1850
rect -3100 1520 3100 1550
rect 3900 4200 10100 4300
rect 10580 4200 10680 5200
rect 3900 2600 10680 4200
rect 3900 1850 10100 2600
rect 3900 1550 4050 1850
rect 9950 1550 10100 1850
rect 3900 1520 10100 1550
rect -3100 1400 10100 1520
rect 10580 1500 10680 2600
rect 10920 1500 11020 7900
rect 10580 1400 11020 1500
rect -7700 300 -6100 1400
rect 1500 1200 5500 1400
rect -4624 880 -4224 881
rect 3300 880 3700 1200
rect -4624 480 3700 880
rect -4624 300 -4224 480
rect -7700 -100 -4224 300
rect -7700 -1200 -6100 -100
rect -12000 -8198 -11060 -4958
rect -10740 -5338 -10420 -5278
rect -10740 -7740 -10698 -5338
rect -10462 -5739 -10420 -5338
rect -10100 -5739 -3900 -1200
rect -1410 -3431 -1010 480
rect -1410 -3711 -1350 -3431
rect -1070 -3711 -1010 -3431
rect -1410 -3771 -1010 -3711
rect -10462 -7339 -3900 -5739
rect -10462 -7740 -10420 -7339
rect -10740 -7800 -10420 -7740
rect -10100 -7350 -3900 -7339
rect -10100 -7650 -9950 -7350
rect -4050 -7650 -3900 -7350
rect -10100 -7800 -3900 -7650
rect -12000 -8300 -11000 -8198
rect -12000 -8900 -11800 -8300
rect -11200 -8900 -11000 -8300
rect -12000 -9000 -11000 -8900
use sky130_fd_sc_hvl__inv_1  sky130_fd_sc_hvl__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1623745244
transform 1 0 -2044 0 -1 -4152
box -66 -43 354 897
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1623745244
transform 1 0 -1756 0 -1 -4152
box -66 -43 834 897
use sky130_fd_pr__pfet_g5v0d10v5_8ATX2D  xm4
timestamp 1623565379
transform 1 0 6000 0 1 -7500
box -1514 -600 1514 600
use sky130_fd_pr__pfet_g5v0d10v5_ZD39PX  xm3
timestamp 1623565379
transform 1 0 6000 0 1 -5700
box -611 -600 611 600
use sky130_fd_sc_hvl__schmittbuf_1  sky130_fd_sc_hvl__schmittbuf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1623745244
transform 1 0 -3100 0 -1 -4152
box -66 -43 1122 897
use sky130_fd_sc_hvl__inv_8  sky130_fd_sc_hvl__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1623745244
transform -1 0 680 0 -1 -4152
box -66 -43 1506 897
use sky130_fd_pr__nfet_g5v0d10v5_7QEKRB  xm2
timestamp 1621758535
transform 1 0 6000 0 1 -1500
box -2351 -588 2351 588
use sky130_fd_pr__nfet_g5v0d10v5_DQEKTK  xm1
timestamp 1621753798
transform 1 0 6000 0 1 -3300
box -3899 -588 3899 588
<< labels >>
flabel metal3 -12000 -5000 -11200 -4600 0 FreeSans 800 0 0 0 iramp
port 1 nsew
flabel metal5 -12000 -9000 -11800 -8200 0 FreeSans 800 0 0 0 vpwr
port 5 nsew
flabel metal3 11200 -5000 12000 -4600 0 FreeSans 800 0 0 0 timeout_int
port 3 nsew
flabel metal4 -10798 320 -10288 800 1 FreeSans 240 0 0 0 vgnd
port 4 n
flabel metal3 11980 -4108 11983 -4008 1 FreeSans 400 0 0 0 rampgen_io
port 2 n
flabel metal3 -2015 -3771 -1989 -3671 1 FreeSans 400 0 0 0 vramp
<< properties >>
string FIXED_BBOX 1158 -4242 10842 -158
<< end >>
