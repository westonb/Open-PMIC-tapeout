magic
tech sky130A
magscale 1 2
timestamp 1623309847
<< nwell >>
rect 1000 -9000 11000 -4600
<< pwell >>
rect 1000 -4400 11000 0
<< mvpsubdiff >>
rect 1066 -78 10934 -66
rect 1066 -238 1300 -78
rect 10700 -238 10934 -78
rect 1066 -250 10934 -238
rect 1066 -300 1250 -250
rect 1066 -4100 1078 -300
rect 1238 -4100 1250 -300
rect 1066 -4150 1250 -4100
rect 10750 -300 10934 -250
rect 10750 -4100 10762 -300
rect 10922 -4100 10934 -300
rect 10750 -4150 10934 -4100
rect 1066 -4162 10934 -4150
rect 1066 -4322 1300 -4162
rect 10700 -4322 10934 -4162
rect 1066 -4334 10934 -4322
<< mvnsubdiff >>
rect 1066 -4678 10934 -4666
rect 1066 -4838 1300 -4678
rect 10700 -4838 10934 -4678
rect 1066 -4850 10934 -4838
rect 1066 -4900 1250 -4850
rect 1066 -8700 1078 -4900
rect 1238 -8700 1250 -4900
rect 1066 -8750 1250 -8700
rect 10750 -4900 10934 -4850
rect 10750 -8700 10762 -4900
rect 10922 -8700 10934 -4900
rect 10750 -8750 10934 -8700
rect 1066 -8762 10934 -8750
rect 1066 -8922 1300 -8762
rect 10700 -8922 10934 -8762
rect 1066 -8934 10934 -8922
<< mvpsubdiffcont >>
rect 1300 -238 10700 -78
rect 1078 -4100 1238 -300
rect 10762 -4100 10922 -300
rect 1300 -4322 10700 -4162
<< mvnsubdiffcont >>
rect 1300 -4838 10700 -4678
rect 1078 -8700 1238 -4900
rect 10762 -8700 10922 -4900
rect 1300 -8922 10700 -8762
<< locali >>
rect 1078 -300 1238 -78
rect 1078 -4322 1238 -4100
rect 10762 -300 10922 -78
rect 10762 -4322 10922 -4100
rect 1078 -4900 1238 -4678
rect 1078 -8922 1238 -8700
rect 10762 -4900 10922 -4678
rect 10762 -8922 10922 -8700
<< viali >>
rect 1238 -238 1300 -78
rect 1300 -238 10700 -78
rect 10700 -238 10762 -78
rect 1078 -3966 1238 -434
rect 10762 -3966 10922 -434
rect 1238 -4322 1300 -4162
rect 1300 -4322 10700 -4162
rect 10700 -4322 10762 -4162
rect 1238 -4838 1300 -4678
rect 1300 -4838 10700 -4678
rect 10700 -4838 10762 -4678
rect 1078 -8566 1238 -5034
rect 10762 -8566 10922 -5034
rect 1238 -8922 1300 -8762
rect 1300 -8922 10700 -8762
rect 10700 -8922 10762 -8762
<< metal1 >>
rect 1072 -78 10928 -72
rect 1072 -238 1238 -78
rect 10762 -238 10928 -78
rect 1072 -244 10928 -238
rect 1072 -434 1244 -244
rect 1072 -3966 1078 -434
rect 1238 -3966 1244 -434
rect 10756 -434 10928 -244
rect 1072 -4156 1244 -3966
rect 1844 -4156 1854 -3856
rect 10146 -4156 10156 -3856
rect 10756 -3966 10762 -434
rect 10922 -3966 10928 -434
rect 10756 -4156 10928 -3966
rect 1072 -4162 10928 -4156
rect 1072 -4322 1238 -4162
rect 10762 -4322 10928 -4162
rect 1072 -4328 10928 -4322
rect 1072 -4678 10928 -4672
rect 1072 -4838 1238 -4678
rect 10762 -4838 10928 -4678
rect 1072 -4844 10928 -4838
rect 1072 -5034 1244 -4844
rect 1072 -8566 1078 -5034
rect 1238 -8566 1244 -5034
rect 1844 -5144 1854 -4844
rect 10146 -5144 10156 -4844
rect 10756 -5034 10928 -4844
rect 1072 -8756 1244 -8566
rect 10756 -8566 10762 -5034
rect 10922 -8566 10928 -5034
rect 10756 -8756 10928 -8566
rect 1072 -8762 10928 -8756
rect 1072 -8922 1238 -8762
rect 10762 -8922 10928 -8762
rect 1072 -8928 10928 -8922
<< via1 >>
rect 1244 -4156 1844 -3856
rect 10156 -4156 10756 -3856
rect 1244 -5144 1844 -4844
rect 10156 -5144 10756 -4844
<< metal2 >>
rect 10237 299 10635 308
rect -8966 -16 -8568 -7
rect -8966 -2706 -8568 -414
rect 10237 -2228 10635 -99
rect 10237 -2721 10651 -2428
rect 11181 -2721 11597 -2720
rect -8966 -3155 -8566 -2906
rect 10237 -3135 11597 -2721
rect -8970 -3545 -8961 -3155
rect -8571 -3545 -8562 -3155
rect -8966 -3550 -8566 -3545
rect 1244 -3856 1844 -3846
rect 1244 -4166 1844 -4156
rect 10156 -3856 10756 -3846
rect 10156 -4166 10756 -4156
rect 11181 -4565 11597 -3135
rect 1244 -4844 1844 -4834
rect 1244 -5154 1844 -5144
rect 10156 -4844 10756 -4834
rect 11181 -4990 11597 -4981
rect 10156 -5154 10756 -5144
<< rmetal2 >>
rect 10237 -2428 10437 -2228
rect -8966 -2906 -8766 -2706
<< via2 >>
rect -8966 -414 -8568 -16
rect 10237 -99 10635 299
rect -8961 -3545 -8571 -3155
rect 1244 -4156 1844 -3856
rect 10156 -4156 10756 -3856
rect 1244 -5144 1844 -4844
rect 10156 -5144 10756 -4844
rect 11181 -4981 11597 -4565
<< metal3 >>
rect 10232 299 10640 304
rect -8971 -16 -8563 -11
rect -9309 -414 -9303 -16
rect -8568 -414 -8563 -16
rect 9488 -99 9494 299
rect 9892 -99 10237 299
rect 10635 -99 10640 299
rect 10232 -104 10640 -99
rect -8971 -419 -8563 -414
rect -8966 -3155 -8566 -3150
rect -8966 -3545 -8961 -3155
rect -8571 -3545 -8566 -3155
rect -8966 -4600 -8566 -3545
rect 1234 -3856 1854 -3851
rect 1234 -4156 1244 -3856
rect 1844 -4156 1854 -3856
rect 1234 -4161 1854 -4156
rect 10146 -3856 10766 -3851
rect 10146 -4156 10156 -3856
rect 10756 -4156 10766 -3856
rect 10146 -4161 10766 -4156
rect -12000 -5000 -8566 -4600
rect 11176 -4565 11602 -4560
rect 1234 -4844 1854 -4839
rect 1234 -5144 1244 -4844
rect 1844 -5144 1854 -4844
rect 1234 -5149 1854 -5144
rect 10146 -4844 10766 -4839
rect 10146 -5144 10156 -4844
rect 10756 -5144 10766 -4844
rect 11176 -4981 11181 -4565
rect 11597 -4600 11602 -4565
rect 11597 -4981 12000 -4600
rect 11176 -4986 12000 -4981
rect 10146 -5149 10766 -5144
rect 11181 -5000 12000 -4986
rect 11181 -5233 11597 -5000
<< via3 >>
rect -9303 -414 -8966 -16
rect -8966 -414 -8905 -16
rect 9494 -99 9892 299
rect 1244 -4156 1844 -3856
rect 10156 -4156 10756 -3856
rect 1244 -5144 1844 -4844
rect 10156 -5144 10756 -4844
<< metal4 >>
rect -12000 8900 12000 9000
rect -12000 8300 -11800 8900
rect -11200 8300 12000 8900
rect -12000 8200 12000 8300
rect -12000 299 12000 800
rect -12000 -16 9494 299
rect -12000 -414 -9303 -16
rect -8905 -99 9494 -16
rect 9892 -99 12000 299
rect -8905 -414 12000 -99
rect -12000 -800 12000 -414
rect 1243 -3856 1845 -3855
rect 1243 -4156 1244 -3856
rect 1844 -4156 1845 -3856
rect 1243 -4157 1845 -4156
rect 10155 -3856 10757 -3855
rect 10155 -4156 10156 -3856
rect 10756 -4156 10757 -3856
rect 10155 -4157 10757 -4156
rect 1243 -4844 1845 -4843
rect 1243 -5144 1244 -4844
rect 1844 -5144 1845 -4844
rect 1243 -5145 1845 -5144
rect 10155 -4844 10757 -4843
rect 10155 -5144 10156 -4844
rect 10756 -5144 10757 -4844
rect 10155 -5145 10757 -5144
rect -12000 -8300 12000 -8200
rect -12000 -8900 -11800 -8300
rect -11200 -8900 12000 -8300
rect -12000 -9000 12000 -8900
<< via4 >>
rect -11800 8300 -11200 8900
rect -11800 -8900 -11200 -8300
<< metal5 >>
rect -12000 8900 -11000 9000
rect -12000 8300 -11800 8900
rect -11200 8300 -11000 8900
rect -12000 -8300 -11000 8300
rect -12000 -8900 -11800 -8300
rect -11200 -8900 -11000 -8300
rect -12000 -9000 -11000 -8900
<< labels >>
flabel metal4 -12000 8200 -12000 9000 3 FreeSans 480 0 0 0 vdd
port 3 e
flabel metal4 -12000 0 -12000 800 3 FreeSans 480 0 0 0 vss
port 4 e
flabel metal3 -12000 -5000 -11200 -4600 0 FreeSans 800 0 0 0 iosc
port 1 nsew
flabel metal3 11200 -5000 12000 -4600 0 FreeSans 800 0 0 0 timeout
port 2 nsew
flabel metal5 -12000 -9000 -11800 -8200 0 FreeSans 800 0 0 0 vdd
port 3 nsew
flabel metal5 -12000 -800 -11800 800 0 FreeSans 800 0 0 0 vss
port 4 nsew
<< properties >>
string FIXED_BBOX 1158 -4242 10842 -158
<< end >>
