magic
tech sky130A
magscale 1 2
timestamp 1624002729
<< metal2 >>
rect -13684 16389 -13584 16398
rect -13884 15795 -13875 15895
rect -13775 15795 -13766 15895
rect -13875 -19421 -13775 15795
rect -13684 -19165 -13584 16289
rect -13496 15095 -13396 15104
rect -13496 -18956 -13396 14995
rect -13139 12797 -12996 12806
rect -13139 12727 -13096 12797
rect -13026 12727 -12996 12797
rect -13139 -18726 -12996 12727
rect -6056 -10643 -5936 -10638
rect -6060 -10753 -6051 -10643
rect -5941 -10753 -5932 -10643
rect -12059 -17937 -11949 -17933
rect -6056 -17937 -5936 -10753
rect -12064 -17942 -11944 -17937
rect -12064 -18052 -12059 -17942
rect -11949 -18052 -11944 -17942
rect -13139 -18869 -12265 -18726
rect -13496 -19056 -12554 -18956
rect -13684 -19265 -12770 -19165
rect -13875 -19521 -12997 -19421
rect -13097 -23750 -12997 -19521
rect -12870 -23585 -12770 -19265
rect -12654 -23415 -12554 -19056
rect -12408 -22918 -12265 -18869
rect -12064 -21147 -11944 -18052
rect -6056 -18066 -5936 -18057
rect -12064 -21276 -11944 -21267
rect -11176 -21355 -11076 -21351
rect -11181 -21360 -11071 -21355
rect -11181 -21460 -11176 -21360
rect -11076 -21460 -11071 -21360
rect -12413 -23051 -12404 -22918
rect -12271 -23051 -12262 -22918
rect -12408 -23055 -12265 -23051
rect -12658 -23505 -12649 -23415
rect -12559 -23505 -12550 -23415
rect -12654 -23510 -12554 -23505
rect -12870 -23675 -12865 -23585
rect -12775 -23675 -12770 -23585
rect -12870 -23680 -12770 -23675
rect -12865 -23684 -12775 -23680
rect -13097 -23859 -12997 -23850
rect -11181 -25273 -11071 -21460
rect -11181 -25392 -11071 -25383
<< via2 >>
rect -13684 16289 -13584 16389
rect -13875 15795 -13775 15895
rect -13496 14995 -13396 15095
rect -13096 12727 -13026 12797
rect -6051 -10753 -5941 -10643
rect -12059 -18052 -11949 -17942
rect -6056 -18057 -5936 -17937
rect -12064 -21267 -11944 -21147
rect -11176 -21460 -11076 -21360
rect -12404 -23051 -12271 -22918
rect -12649 -23505 -12559 -23415
rect -12865 -23675 -12775 -23585
rect -13097 -23850 -12997 -23750
rect -11181 -25383 -11071 -25273
<< metal3 >>
rect -13689 16389 -13579 16394
rect -13689 16289 -13684 16389
rect -13584 16289 -10494 16389
rect -13689 16284 -13579 16289
rect -13880 15895 -13770 15900
rect -13880 15795 -13875 15895
rect -13775 15795 -10486 15895
rect -13880 15790 -13770 15795
rect -18203 15363 -10455 15439
rect -13501 15095 -13391 15100
rect -10514 15095 -10314 15122
rect -13501 14995 -13496 15095
rect -13396 14995 -10314 15095
rect -13501 14990 -13391 14995
rect -18210 14799 -10429 14879
rect 11664 14238 11825 14326
rect 11684 13474 11792 13534
rect -13101 12797 -10416 12802
rect -13101 12727 -13096 12797
rect -13026 12727 -10416 12797
rect -13101 12722 -10416 12727
rect 11668 9916 11786 9988
rect -10564 7772 -9918 8172
rect -10564 -1321 -10164 7772
rect 11286 -1232 12079 -992
rect 11417 -1540 12083 -1440
rect 11431 -1864 12083 -1764
rect -17951 -7724 -11546 -7464
rect -6370 -10643 -5936 -10638
rect -6370 -10753 -6051 -10643
rect -5941 -10753 -5936 -10643
rect -6370 -10758 -5936 -10753
rect -6061 -17937 -5931 -17932
rect -12064 -17942 -6056 -17937
rect -12064 -18052 -12059 -17942
rect -11949 -18052 -6056 -17942
rect -12064 -18057 -6056 -18052
rect -5936 -18057 -5931 -17937
rect -6061 -18062 -5931 -18057
rect -12069 -21147 -11939 -21142
rect -13143 -21267 -12064 -21147
rect -11944 -21267 -11939 -21147
rect -12069 -21272 -11939 -21267
rect -13199 -21360 -11071 -21355
rect -13199 -21460 -11176 -21360
rect -11076 -21460 -11071 -21360
rect -13199 -21465 -11071 -21460
rect -18154 -22459 -11436 -22359
rect -18152 -22704 -11445 -22604
rect -10049 -22610 4945 -22410
rect -10049 -22885 -9849 -22610
rect -18173 -22918 -9849 -22885
rect -18173 -23051 -12404 -22918
rect -12271 -23051 -9849 -22918
rect -18173 -23085 -9849 -23051
rect -12654 -23415 -12554 -23410
rect -12654 -23505 -12649 -23415
rect -12559 -23505 -12554 -23415
rect -12654 -23510 -12554 -23505
rect -12870 -23585 -12589 -23580
rect -12870 -23675 -12865 -23585
rect -12775 -23675 -12589 -23585
rect -12870 -23680 -12589 -23675
rect -13102 -23750 -12992 -23745
rect -13102 -23850 -13097 -23750
rect -12997 -23850 -12992 -23750
rect -13102 -23855 -12992 -23850
rect -11186 -25273 -11066 -25268
rect -18100 -25480 -17328 -25280
rect -11186 -25383 -11181 -25273
rect -11071 -25383 -11066 -25273
rect -11186 -25388 -11066 -25383
<< metal4 >>
rect -19000 18741 13000 18800
rect -19000 17260 12120 18741
rect 12900 17260 13000 18741
rect -19000 17200 13000 17260
rect -19000 9741 13000 9800
rect -19000 8260 -18940 9741
rect -18160 8260 13000 9741
rect -19000 8200 13000 8260
rect -19000 741 13000 800
rect -19000 -740 12120 741
rect 12900 -740 13000 741
rect -19000 -800 13000 -740
rect -19000 -8259 13000 -8200
rect -19000 -9740 -18940 -8259
rect -18160 -9740 13000 -8259
rect -19000 -9800 13000 -9740
rect -19000 -17259 13000 -17200
rect -19000 -18740 12120 -17259
rect 12900 -18740 13000 -17259
rect -19000 -18800 13000 -18740
rect -19000 -26259 13000 -26200
rect -19000 -27740 -18940 -26259
rect -18160 -27740 13000 -26259
rect -19000 -27800 13000 -27740
<< via4 >>
rect 12120 17260 12900 18741
rect -18940 8260 -18160 9741
rect 12120 -740 12900 741
rect -18940 -9740 -18160 -8259
rect 12120 -18740 12900 -17259
rect -18940 -27740 -18160 -26259
<< metal5 >>
rect -19000 9741 -18000 18800
rect -19000 8260 -18940 9741
rect -18160 8260 -18000 9741
rect -19000 -8259 -18000 8260
rect -19000 -9740 -18940 -8259
rect -18160 -9740 -18000 -8259
rect -19000 -26259 -18000 -9740
rect -19000 -27740 -18940 -26259
rect -18160 -27740 -18000 -26259
rect -19000 -27800 -18000 -27740
rect 12000 18741 13000 18800
rect 12000 17260 12120 18741
rect 12900 17260 13000 18741
rect 12000 741 13000 17260
rect 12000 -740 12120 741
rect 12900 -740 13000 741
rect 12000 -17259 13000 -740
rect 12000 -18740 12120 -17259
rect 12900 -18740 13000 -17259
rect 12000 -27800 13000 -18740
use modulator  modulator_0
timestamp 1624002729
transform 1 0 0 0 -1 9000
box -12000 -9000 12000 9000
use bias_distribution  bias_distribution_0
timestamp 1624002729
transform 1 0 -15000 0 1 -22500
box -3000 -4500 3000 4500
use current_sense  current_sense_0
timestamp 1624002729
transform -1 0 0 0 1 -9000
box -12000 -9000 12000 9000
use folded_cascode_p_in  folded_cascode_p_in_0
timestamp 1624002729
transform 1 0 -3000 0 1 -22500
box -9000 -4500 15000 4500
<< labels >>
flabel metal3 -18154 -22459 -18152 -22359 3 FreeSans 400 0 0 0 vref
port 14 e
flabel metal3 -18152 -22704 -18150 -22604 3 FreeSans 400 0 0 0 vfb
port 13 e
flabel metal3 -18100 -25480 -18097 -25280 1 FreeSans 400 0 0 0 ibias
port 2 n
flabel metal3 11823 14238 11825 14326 1 FreeSans 400 0 0 0 overcurrent
port 6 n
flabel metal3 11791 13474 11792 13534 1 FreeSans 400 0 0 0 cycle_end
port 1 n
flabel metal3 -18173 -23085 -18168 -22885 1 FreeSans 400 0 0 0 vcomp
port 11 n
flabel metal3 -18203 15363 -18200 15439 1 FreeSans 400 0 0 0 islope
port 5 n
flabel metal3 -18210 14799 -18207 14879 3 FreeSans 400 0 0 0 ioc
port 4 e
flabel metal3 11784 9916 11786 9988 1 FreeSans 400 0 0 0 timeout
port 10 n
flabel metal3 -17951 -7724 -17946 -7464 1 FreeSans 400 0 0 0 imon
port 3 n
flabel metal3 12076 -1232 12079 -992 1 FreeSans 400 0 0 0 sense_fet
port 7 n
flabel metal3 12081 -1540 12083 -1440 7 FreeSans 400 0 0 0 sense_fet_kelvin
port 8 w
flabel metal3 12081 -1864 12083 -1764 7 FreeSans 400 0 0 0 sw_node
port 9 w
flabel metal4 -19000 -27800 -18997 -26200 0 FreeSans 400 0 0 0 vss
port 15 nsew
flabel metal4 -19000 -18800 -18997 -17200 0 FreeSans 400 0 0 0 vdd
port 12 nsew
<< end >>
