magic
tech sky130A
magscale 1 2
timestamp 1624002729
<< error_p >>
rect -1319 -500 -1261 500
rect -1061 -500 -1003 500
rect -803 -500 -745 500
rect -545 -500 -487 500
rect -287 -500 -229 500
rect -29 -500 29 500
rect 229 -500 287 500
rect 487 -500 545 500
rect 745 -500 803 500
rect 1003 -500 1061 500
rect 1261 -500 1319 500
<< mvnmos >>
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
<< mvndiff >>
rect -1319 488 -1261 500
rect -1319 -488 -1307 488
rect -1273 -488 -1261 488
rect -1319 -500 -1261 -488
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
rect 1261 488 1319 500
rect 1261 -488 1273 488
rect 1307 -488 1319 488
rect 1261 -500 1319 -488
<< mvndiffc >>
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
<< poly >>
rect -1227 572 -1095 588
rect -1227 555 -1211 572
rect -1261 538 -1211 555
rect -1111 555 -1095 572
rect -969 572 -837 588
rect -969 555 -953 572
rect -1111 538 -1061 555
rect -1261 500 -1061 538
rect -1003 538 -953 555
rect -853 555 -837 572
rect -711 572 -579 588
rect -711 555 -695 572
rect -853 538 -803 555
rect -1003 500 -803 538
rect -745 538 -695 555
rect -595 555 -579 572
rect -453 572 -321 588
rect -453 555 -437 572
rect -595 538 -545 555
rect -745 500 -545 538
rect -487 538 -437 555
rect -337 555 -321 572
rect -195 572 -63 588
rect -195 555 -179 572
rect -337 538 -287 555
rect -487 500 -287 538
rect -229 538 -179 555
rect -79 555 -63 572
rect 63 572 195 588
rect 63 555 79 572
rect -79 538 -29 555
rect -229 500 -29 538
rect 29 538 79 555
rect 179 555 195 572
rect 321 572 453 588
rect 321 555 337 572
rect 179 538 229 555
rect 29 500 229 538
rect 287 538 337 555
rect 437 555 453 572
rect 579 572 711 588
rect 579 555 595 572
rect 437 538 487 555
rect 287 500 487 538
rect 545 538 595 555
rect 695 555 711 572
rect 837 572 969 588
rect 837 555 853 572
rect 695 538 745 555
rect 545 500 745 538
rect 803 538 853 555
rect 953 555 969 572
rect 1095 572 1227 588
rect 1095 555 1111 572
rect 953 538 1003 555
rect 803 500 1003 538
rect 1061 538 1111 555
rect 1211 555 1227 572
rect 1211 538 1261 555
rect 1061 500 1261 538
rect -1261 -538 -1061 -500
rect -1261 -555 -1211 -538
rect -1227 -572 -1211 -555
rect -1111 -555 -1061 -538
rect -1003 -538 -803 -500
rect -1003 -555 -953 -538
rect -1111 -572 -1095 -555
rect -1227 -588 -1095 -572
rect -969 -572 -953 -555
rect -853 -555 -803 -538
rect -745 -538 -545 -500
rect -745 -555 -695 -538
rect -853 -572 -837 -555
rect -969 -588 -837 -572
rect -711 -572 -695 -555
rect -595 -555 -545 -538
rect -487 -538 -287 -500
rect -487 -555 -437 -538
rect -595 -572 -579 -555
rect -711 -588 -579 -572
rect -453 -572 -437 -555
rect -337 -555 -287 -538
rect -229 -538 -29 -500
rect -229 -555 -179 -538
rect -337 -572 -321 -555
rect -453 -588 -321 -572
rect -195 -572 -179 -555
rect -79 -555 -29 -538
rect 29 -538 229 -500
rect 29 -555 79 -538
rect -79 -572 -63 -555
rect -195 -588 -63 -572
rect 63 -572 79 -555
rect 179 -555 229 -538
rect 287 -538 487 -500
rect 287 -555 337 -538
rect 179 -572 195 -555
rect 63 -588 195 -572
rect 321 -572 337 -555
rect 437 -555 487 -538
rect 545 -538 745 -500
rect 545 -555 595 -538
rect 437 -572 453 -555
rect 321 -588 453 -572
rect 579 -572 595 -555
rect 695 -555 745 -538
rect 803 -538 1003 -500
rect 803 -555 853 -538
rect 695 -572 711 -555
rect 579 -588 711 -572
rect 837 -572 853 -555
rect 953 -555 1003 -538
rect 1061 -538 1261 -500
rect 1061 -555 1111 -538
rect 953 -572 969 -555
rect 837 -588 969 -572
rect 1095 -572 1111 -555
rect 1211 -555 1261 -538
rect 1211 -572 1227 -555
rect 1095 -588 1227 -572
<< polycont >>
rect -1211 538 -1111 572
rect -953 538 -853 572
rect -695 538 -595 572
rect -437 538 -337 572
rect -179 538 -79 572
rect 79 538 179 572
rect 337 538 437 572
rect 595 538 695 572
rect 853 538 953 572
rect 1111 538 1211 572
rect -1211 -572 -1111 -538
rect -953 -572 -853 -538
rect -695 -572 -595 -538
rect -437 -572 -337 -538
rect -179 -572 -79 -538
rect 79 -572 179 -538
rect 337 -572 437 -538
rect 595 -572 695 -538
rect 853 -572 953 -538
rect 1111 -572 1211 -538
<< locali >>
rect -1227 538 -1211 572
rect -1111 538 -1095 572
rect -969 538 -953 572
rect -853 538 -837 572
rect -711 538 -695 572
rect -595 538 -579 572
rect -453 538 -437 572
rect -337 538 -321 572
rect -195 538 -179 572
rect -79 538 -63 572
rect 63 538 79 572
rect 179 538 195 572
rect 321 538 337 572
rect 437 538 453 572
rect 579 538 595 572
rect 695 538 711 572
rect 837 538 853 572
rect 953 538 969 572
rect 1095 538 1111 572
rect 1211 538 1227 572
rect -1307 488 -1273 504
rect -1307 -504 -1273 -488
rect -1049 488 -1015 504
rect -1049 -504 -1015 -488
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -504 1049 -488
rect 1273 488 1307 504
rect 1273 -504 1307 -488
rect -1227 -572 -1211 -538
rect -1111 -572 -1095 -538
rect -969 -572 -953 -538
rect -853 -572 -837 -538
rect -711 -572 -695 -538
rect -595 -572 -579 -538
rect -453 -572 -437 -538
rect -337 -572 -321 -538
rect -195 -572 -179 -538
rect -79 -572 -63 -538
rect 63 -572 79 -538
rect 179 -572 195 -538
rect 321 -572 337 -538
rect 437 -572 453 -538
rect 579 -572 595 -538
rect 695 -572 711 -538
rect 837 -572 853 -538
rect 953 -572 969 -538
rect 1095 -572 1111 -538
rect 1211 -572 1227 -538
<< viali >>
rect -1195 538 -1127 572
rect -937 538 -869 572
rect -679 538 -611 572
rect -421 538 -353 572
rect -163 538 -95 572
rect 95 538 163 572
rect 353 538 421 572
rect 611 538 679 572
rect 869 538 937 572
rect 1127 538 1195 572
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect -1195 -572 -1127 -538
rect -937 -572 -869 -538
rect -679 -572 -611 -538
rect -421 -572 -353 -538
rect -163 -572 -95 -538
rect 95 -572 163 -538
rect 353 -572 421 -538
rect 611 -572 679 -538
rect 869 -572 937 -538
rect 1127 -572 1195 -538
<< metal1 >>
rect -1207 572 -1115 578
rect -1207 538 -1195 572
rect -1127 538 -1115 572
rect -1207 532 -1115 538
rect -949 572 -857 578
rect -949 538 -937 572
rect -869 538 -857 572
rect -949 532 -857 538
rect -691 572 -599 578
rect -691 538 -679 572
rect -611 538 -599 572
rect -691 532 -599 538
rect -433 572 -341 578
rect -433 538 -421 572
rect -353 538 -341 572
rect -433 532 -341 538
rect -175 572 -83 578
rect -175 538 -163 572
rect -95 538 -83 572
rect -175 532 -83 538
rect 83 572 175 578
rect 83 538 95 572
rect 163 538 175 572
rect 83 532 175 538
rect 341 572 433 578
rect 341 538 353 572
rect 421 538 433 572
rect 341 532 433 538
rect 599 572 691 578
rect 599 538 611 572
rect 679 538 691 572
rect 599 532 691 538
rect 857 572 949 578
rect 857 538 869 572
rect 937 538 949 572
rect 857 532 949 538
rect 1115 572 1207 578
rect 1115 538 1127 572
rect 1195 538 1207 572
rect 1115 532 1207 538
rect -1313 488 -1267 500
rect -1313 -488 -1307 488
rect -1273 -488 -1267 488
rect -1313 -500 -1267 -488
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect 1267 488 1313 500
rect 1267 -488 1273 488
rect 1307 -488 1313 488
rect 1267 -500 1313 -488
rect -1207 -538 -1115 -532
rect -1207 -572 -1195 -538
rect -1127 -572 -1115 -538
rect -1207 -578 -1115 -572
rect -949 -538 -857 -532
rect -949 -572 -937 -538
rect -869 -572 -857 -538
rect -949 -578 -857 -572
rect -691 -538 -599 -532
rect -691 -572 -679 -538
rect -611 -572 -599 -538
rect -691 -578 -599 -572
rect -433 -538 -341 -532
rect -433 -572 -421 -538
rect -353 -572 -341 -538
rect -433 -578 -341 -572
rect -175 -538 -83 -532
rect -175 -572 -163 -538
rect -95 -572 -83 -538
rect -175 -578 -83 -572
rect 83 -538 175 -532
rect 83 -572 95 -538
rect 163 -572 175 -538
rect 83 -578 175 -572
rect 341 -538 433 -532
rect 341 -572 353 -538
rect 421 -572 433 -538
rect 341 -578 433 -572
rect 599 -538 691 -532
rect 599 -572 611 -538
rect 679 -572 691 -538
rect 599 -578 691 -572
rect 857 -538 949 -532
rect 857 -572 869 -538
rect 937 -572 949 -538
rect 857 -578 949 -572
rect 1115 -538 1207 -532
rect 1115 -572 1127 -538
rect 1195 -572 1207 -538
rect 1115 -578 1207 -572
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string parameters w 5 l 1 m 1 nf 10 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
