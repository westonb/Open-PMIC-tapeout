magic
tech sky130A
magscale 1 2
timestamp 1624002729
<< error_p >>
rect -4645 566 4645 600
rect -4675 -566 4675 566
rect -4645 -600 4645 -566
<< nwell >>
rect -4645 -600 4645 600
<< mvpmos >>
rect -4551 -500 -4151 500
rect -4093 -500 -3693 500
rect -3635 -500 -3235 500
rect -3177 -500 -2777 500
rect -2719 -500 -2319 500
rect -2261 -500 -1861 500
rect -1803 -500 -1403 500
rect -1345 -500 -945 500
rect -887 -500 -487 500
rect -429 -500 -29 500
rect 29 -500 429 500
rect 487 -500 887 500
rect 945 -500 1345 500
rect 1403 -500 1803 500
rect 1861 -500 2261 500
rect 2319 -500 2719 500
rect 2777 -500 3177 500
rect 3235 -500 3635 500
rect 3693 -500 4093 500
rect 4151 -500 4551 500
<< mvpdiff >>
rect -4609 488 -4551 500
rect -4609 -488 -4597 488
rect -4563 -488 -4551 488
rect -4609 -500 -4551 -488
rect -4151 488 -4093 500
rect -4151 -488 -4139 488
rect -4105 -488 -4093 488
rect -4151 -500 -4093 -488
rect -3693 488 -3635 500
rect -3693 -488 -3681 488
rect -3647 -488 -3635 488
rect -3693 -500 -3635 -488
rect -3235 488 -3177 500
rect -3235 -488 -3223 488
rect -3189 -488 -3177 488
rect -3235 -500 -3177 -488
rect -2777 488 -2719 500
rect -2777 -488 -2765 488
rect -2731 -488 -2719 488
rect -2777 -500 -2719 -488
rect -2319 488 -2261 500
rect -2319 -488 -2307 488
rect -2273 -488 -2261 488
rect -2319 -500 -2261 -488
rect -1861 488 -1803 500
rect -1861 -488 -1849 488
rect -1815 -488 -1803 488
rect -1861 -500 -1803 -488
rect -1403 488 -1345 500
rect -1403 -488 -1391 488
rect -1357 -488 -1345 488
rect -1403 -500 -1345 -488
rect -945 488 -887 500
rect -945 -488 -933 488
rect -899 -488 -887 488
rect -945 -500 -887 -488
rect -487 488 -429 500
rect -487 -488 -475 488
rect -441 -488 -429 488
rect -487 -500 -429 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 429 488 487 500
rect 429 -488 441 488
rect 475 -488 487 488
rect 429 -500 487 -488
rect 887 488 945 500
rect 887 -488 899 488
rect 933 -488 945 488
rect 887 -500 945 -488
rect 1345 488 1403 500
rect 1345 -488 1357 488
rect 1391 -488 1403 488
rect 1345 -500 1403 -488
rect 1803 488 1861 500
rect 1803 -488 1815 488
rect 1849 -488 1861 488
rect 1803 -500 1861 -488
rect 2261 488 2319 500
rect 2261 -488 2273 488
rect 2307 -488 2319 488
rect 2261 -500 2319 -488
rect 2719 488 2777 500
rect 2719 -488 2731 488
rect 2765 -488 2777 488
rect 2719 -500 2777 -488
rect 3177 488 3235 500
rect 3177 -488 3189 488
rect 3223 -488 3235 488
rect 3177 -500 3235 -488
rect 3635 488 3693 500
rect 3635 -488 3647 488
rect 3681 -488 3693 488
rect 3635 -500 3693 -488
rect 4093 488 4151 500
rect 4093 -488 4105 488
rect 4139 -488 4151 488
rect 4093 -500 4151 -488
rect 4551 488 4609 500
rect 4551 -488 4563 488
rect 4597 -488 4609 488
rect 4551 -500 4609 -488
<< mvpdiffc >>
rect -4597 -488 -4563 488
rect -4139 -488 -4105 488
rect -3681 -488 -3647 488
rect -3223 -488 -3189 488
rect -2765 -488 -2731 488
rect -2307 -488 -2273 488
rect -1849 -488 -1815 488
rect -1391 -488 -1357 488
rect -933 -488 -899 488
rect -475 -488 -441 488
rect -17 -488 17 488
rect 441 -488 475 488
rect 899 -488 933 488
rect 1357 -488 1391 488
rect 1815 -488 1849 488
rect 2273 -488 2307 488
rect 2731 -488 2765 488
rect 3189 -488 3223 488
rect 3647 -488 3681 488
rect 4105 -488 4139 488
rect 4563 -488 4597 488
<< poly >>
rect -4477 581 -4225 597
rect -4477 564 -4461 581
rect -4551 547 -4461 564
rect -4241 564 -4225 581
rect -4019 581 -3767 597
rect -4019 564 -4003 581
rect -4241 547 -4151 564
rect -4551 500 -4151 547
rect -4093 547 -4003 564
rect -3783 564 -3767 581
rect -3561 581 -3309 597
rect -3561 564 -3545 581
rect -3783 547 -3693 564
rect -4093 500 -3693 547
rect -3635 547 -3545 564
rect -3325 564 -3309 581
rect -3103 581 -2851 597
rect -3103 564 -3087 581
rect -3325 547 -3235 564
rect -3635 500 -3235 547
rect -3177 547 -3087 564
rect -2867 564 -2851 581
rect -2645 581 -2393 597
rect -2645 564 -2629 581
rect -2867 547 -2777 564
rect -3177 500 -2777 547
rect -2719 547 -2629 564
rect -2409 564 -2393 581
rect -2187 581 -1935 597
rect -2187 564 -2171 581
rect -2409 547 -2319 564
rect -2719 500 -2319 547
rect -2261 547 -2171 564
rect -1951 564 -1935 581
rect -1729 581 -1477 597
rect -1729 564 -1713 581
rect -1951 547 -1861 564
rect -2261 500 -1861 547
rect -1803 547 -1713 564
rect -1493 564 -1477 581
rect -1271 581 -1019 597
rect -1271 564 -1255 581
rect -1493 547 -1403 564
rect -1803 500 -1403 547
rect -1345 547 -1255 564
rect -1035 564 -1019 581
rect -813 581 -561 597
rect -813 564 -797 581
rect -1035 547 -945 564
rect -1345 500 -945 547
rect -887 547 -797 564
rect -577 564 -561 581
rect -355 581 -103 597
rect -355 564 -339 581
rect -577 547 -487 564
rect -887 500 -487 547
rect -429 547 -339 564
rect -119 564 -103 581
rect 103 581 355 597
rect 103 564 119 581
rect -119 547 -29 564
rect -429 500 -29 547
rect 29 547 119 564
rect 339 564 355 581
rect 561 581 813 597
rect 561 564 577 581
rect 339 547 429 564
rect 29 500 429 547
rect 487 547 577 564
rect 797 564 813 581
rect 1019 581 1271 597
rect 1019 564 1035 581
rect 797 547 887 564
rect 487 500 887 547
rect 945 547 1035 564
rect 1255 564 1271 581
rect 1477 581 1729 597
rect 1477 564 1493 581
rect 1255 547 1345 564
rect 945 500 1345 547
rect 1403 547 1493 564
rect 1713 564 1729 581
rect 1935 581 2187 597
rect 1935 564 1951 581
rect 1713 547 1803 564
rect 1403 500 1803 547
rect 1861 547 1951 564
rect 2171 564 2187 581
rect 2393 581 2645 597
rect 2393 564 2409 581
rect 2171 547 2261 564
rect 1861 500 2261 547
rect 2319 547 2409 564
rect 2629 564 2645 581
rect 2851 581 3103 597
rect 2851 564 2867 581
rect 2629 547 2719 564
rect 2319 500 2719 547
rect 2777 547 2867 564
rect 3087 564 3103 581
rect 3309 581 3561 597
rect 3309 564 3325 581
rect 3087 547 3177 564
rect 2777 500 3177 547
rect 3235 547 3325 564
rect 3545 564 3561 581
rect 3767 581 4019 597
rect 3767 564 3783 581
rect 3545 547 3635 564
rect 3235 500 3635 547
rect 3693 547 3783 564
rect 4003 564 4019 581
rect 4225 581 4477 597
rect 4225 564 4241 581
rect 4003 547 4093 564
rect 3693 500 4093 547
rect 4151 547 4241 564
rect 4461 564 4477 581
rect 4461 547 4551 564
rect 4151 500 4551 547
rect -4551 -547 -4151 -500
rect -4551 -564 -4461 -547
rect -4477 -581 -4461 -564
rect -4241 -564 -4151 -547
rect -4093 -547 -3693 -500
rect -4093 -564 -4003 -547
rect -4241 -581 -4225 -564
rect -4477 -597 -4225 -581
rect -4019 -581 -4003 -564
rect -3783 -564 -3693 -547
rect -3635 -547 -3235 -500
rect -3635 -564 -3545 -547
rect -3783 -581 -3767 -564
rect -4019 -597 -3767 -581
rect -3561 -581 -3545 -564
rect -3325 -564 -3235 -547
rect -3177 -547 -2777 -500
rect -3177 -564 -3087 -547
rect -3325 -581 -3309 -564
rect -3561 -597 -3309 -581
rect -3103 -581 -3087 -564
rect -2867 -564 -2777 -547
rect -2719 -547 -2319 -500
rect -2719 -564 -2629 -547
rect -2867 -581 -2851 -564
rect -3103 -597 -2851 -581
rect -2645 -581 -2629 -564
rect -2409 -564 -2319 -547
rect -2261 -547 -1861 -500
rect -2261 -564 -2171 -547
rect -2409 -581 -2393 -564
rect -2645 -597 -2393 -581
rect -2187 -581 -2171 -564
rect -1951 -564 -1861 -547
rect -1803 -547 -1403 -500
rect -1803 -564 -1713 -547
rect -1951 -581 -1935 -564
rect -2187 -597 -1935 -581
rect -1729 -581 -1713 -564
rect -1493 -564 -1403 -547
rect -1345 -547 -945 -500
rect -1345 -564 -1255 -547
rect -1493 -581 -1477 -564
rect -1729 -597 -1477 -581
rect -1271 -581 -1255 -564
rect -1035 -564 -945 -547
rect -887 -547 -487 -500
rect -887 -564 -797 -547
rect -1035 -581 -1019 -564
rect -1271 -597 -1019 -581
rect -813 -581 -797 -564
rect -577 -564 -487 -547
rect -429 -547 -29 -500
rect -429 -564 -339 -547
rect -577 -581 -561 -564
rect -813 -597 -561 -581
rect -355 -581 -339 -564
rect -119 -564 -29 -547
rect 29 -547 429 -500
rect 29 -564 119 -547
rect -119 -581 -103 -564
rect -355 -597 -103 -581
rect 103 -581 119 -564
rect 339 -564 429 -547
rect 487 -547 887 -500
rect 487 -564 577 -547
rect 339 -581 355 -564
rect 103 -597 355 -581
rect 561 -581 577 -564
rect 797 -564 887 -547
rect 945 -547 1345 -500
rect 945 -564 1035 -547
rect 797 -581 813 -564
rect 561 -597 813 -581
rect 1019 -581 1035 -564
rect 1255 -564 1345 -547
rect 1403 -547 1803 -500
rect 1403 -564 1493 -547
rect 1255 -581 1271 -564
rect 1019 -597 1271 -581
rect 1477 -581 1493 -564
rect 1713 -564 1803 -547
rect 1861 -547 2261 -500
rect 1861 -564 1951 -547
rect 1713 -581 1729 -564
rect 1477 -597 1729 -581
rect 1935 -581 1951 -564
rect 2171 -564 2261 -547
rect 2319 -547 2719 -500
rect 2319 -564 2409 -547
rect 2171 -581 2187 -564
rect 1935 -597 2187 -581
rect 2393 -581 2409 -564
rect 2629 -564 2719 -547
rect 2777 -547 3177 -500
rect 2777 -564 2867 -547
rect 2629 -581 2645 -564
rect 2393 -597 2645 -581
rect 2851 -581 2867 -564
rect 3087 -564 3177 -547
rect 3235 -547 3635 -500
rect 3235 -564 3325 -547
rect 3087 -581 3103 -564
rect 2851 -597 3103 -581
rect 3309 -581 3325 -564
rect 3545 -564 3635 -547
rect 3693 -547 4093 -500
rect 3693 -564 3783 -547
rect 3545 -581 3561 -564
rect 3309 -597 3561 -581
rect 3767 -581 3783 -564
rect 4003 -564 4093 -547
rect 4151 -547 4551 -500
rect 4151 -564 4241 -547
rect 4003 -581 4019 -564
rect 3767 -597 4019 -581
rect 4225 -581 4241 -564
rect 4461 -564 4551 -547
rect 4461 -581 4477 -564
rect 4225 -597 4477 -581
<< polycont >>
rect -4461 547 -4241 581
rect -4003 547 -3783 581
rect -3545 547 -3325 581
rect -3087 547 -2867 581
rect -2629 547 -2409 581
rect -2171 547 -1951 581
rect -1713 547 -1493 581
rect -1255 547 -1035 581
rect -797 547 -577 581
rect -339 547 -119 581
rect 119 547 339 581
rect 577 547 797 581
rect 1035 547 1255 581
rect 1493 547 1713 581
rect 1951 547 2171 581
rect 2409 547 2629 581
rect 2867 547 3087 581
rect 3325 547 3545 581
rect 3783 547 4003 581
rect 4241 547 4461 581
rect -4461 -581 -4241 -547
rect -4003 -581 -3783 -547
rect -3545 -581 -3325 -547
rect -3087 -581 -2867 -547
rect -2629 -581 -2409 -547
rect -2171 -581 -1951 -547
rect -1713 -581 -1493 -547
rect -1255 -581 -1035 -547
rect -797 -581 -577 -547
rect -339 -581 -119 -547
rect 119 -581 339 -547
rect 577 -581 797 -547
rect 1035 -581 1255 -547
rect 1493 -581 1713 -547
rect 1951 -581 2171 -547
rect 2409 -581 2629 -547
rect 2867 -581 3087 -547
rect 3325 -581 3545 -547
rect 3783 -581 4003 -547
rect 4241 -581 4461 -547
<< locali >>
rect -4477 547 -4461 581
rect -4241 547 -4225 581
rect -4019 547 -4003 581
rect -3783 547 -3767 581
rect -3561 547 -3545 581
rect -3325 547 -3309 581
rect -3103 547 -3087 581
rect -2867 547 -2851 581
rect -2645 547 -2629 581
rect -2409 547 -2393 581
rect -2187 547 -2171 581
rect -1951 547 -1935 581
rect -1729 547 -1713 581
rect -1493 547 -1477 581
rect -1271 547 -1255 581
rect -1035 547 -1019 581
rect -813 547 -797 581
rect -577 547 -561 581
rect -355 547 -339 581
rect -119 547 -103 581
rect 103 547 119 581
rect 339 547 355 581
rect 561 547 577 581
rect 797 547 813 581
rect 1019 547 1035 581
rect 1255 547 1271 581
rect 1477 547 1493 581
rect 1713 547 1729 581
rect 1935 547 1951 581
rect 2171 547 2187 581
rect 2393 547 2409 581
rect 2629 547 2645 581
rect 2851 547 2867 581
rect 3087 547 3103 581
rect 3309 547 3325 581
rect 3545 547 3561 581
rect 3767 547 3783 581
rect 4003 547 4019 581
rect 4225 547 4241 581
rect 4461 547 4477 581
rect -4597 488 -4563 504
rect -4597 -504 -4563 -488
rect -4139 488 -4105 504
rect -4139 -504 -4105 -488
rect -3681 488 -3647 504
rect -3681 -504 -3647 -488
rect -3223 488 -3189 504
rect -3223 -504 -3189 -488
rect -2765 488 -2731 504
rect -2765 -504 -2731 -488
rect -2307 488 -2273 504
rect -2307 -504 -2273 -488
rect -1849 488 -1815 504
rect -1849 -504 -1815 -488
rect -1391 488 -1357 504
rect -1391 -504 -1357 -488
rect -933 488 -899 504
rect -933 -504 -899 -488
rect -475 488 -441 504
rect -475 -504 -441 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 441 488 475 504
rect 441 -504 475 -488
rect 899 488 933 504
rect 899 -504 933 -488
rect 1357 488 1391 504
rect 1357 -504 1391 -488
rect 1815 488 1849 504
rect 1815 -504 1849 -488
rect 2273 488 2307 504
rect 2273 -504 2307 -488
rect 2731 488 2765 504
rect 2731 -504 2765 -488
rect 3189 488 3223 504
rect 3189 -504 3223 -488
rect 3647 488 3681 504
rect 3647 -504 3681 -488
rect 4105 488 4139 504
rect 4105 -504 4139 -488
rect 4563 488 4597 504
rect 4563 -504 4597 -488
rect -4477 -581 -4461 -547
rect -4241 -581 -4225 -547
rect -4019 -581 -4003 -547
rect -3783 -581 -3767 -547
rect -3561 -581 -3545 -547
rect -3325 -581 -3309 -547
rect -3103 -581 -3087 -547
rect -2867 -581 -2851 -547
rect -2645 -581 -2629 -547
rect -2409 -581 -2393 -547
rect -2187 -581 -2171 -547
rect -1951 -581 -1935 -547
rect -1729 -581 -1713 -547
rect -1493 -581 -1477 -547
rect -1271 -581 -1255 -547
rect -1035 -581 -1019 -547
rect -813 -581 -797 -547
rect -577 -581 -561 -547
rect -355 -581 -339 -547
rect -119 -581 -103 -547
rect 103 -581 119 -547
rect 339 -581 355 -547
rect 561 -581 577 -547
rect 797 -581 813 -547
rect 1019 -581 1035 -547
rect 1255 -581 1271 -547
rect 1477 -581 1493 -547
rect 1713 -581 1729 -547
rect 1935 -581 1951 -547
rect 2171 -581 2187 -547
rect 2393 -581 2409 -547
rect 2629 -581 2645 -547
rect 2851 -581 2867 -547
rect 3087 -581 3103 -547
rect 3309 -581 3325 -547
rect 3545 -581 3561 -547
rect 3767 -581 3783 -547
rect 4003 -581 4019 -547
rect 4225 -581 4241 -547
rect 4461 -581 4477 -547
<< viali >>
rect -4425 547 -4277 581
rect -3967 547 -3819 581
rect -3509 547 -3361 581
rect -3051 547 -2903 581
rect -2593 547 -2445 581
rect -2135 547 -1987 581
rect -1677 547 -1529 581
rect -1219 547 -1071 581
rect -761 547 -613 581
rect -303 547 -155 581
rect 155 547 303 581
rect 613 547 761 581
rect 1071 547 1219 581
rect 1529 547 1677 581
rect 1987 547 2135 581
rect 2445 547 2593 581
rect 2903 547 3051 581
rect 3361 547 3509 581
rect 3819 547 3967 581
rect 4277 547 4425 581
rect -4597 -488 -4563 488
rect -4139 -488 -4105 488
rect -3681 -488 -3647 488
rect -3223 -488 -3189 488
rect -2765 -488 -2731 488
rect -2307 -488 -2273 488
rect -1849 -488 -1815 488
rect -1391 -488 -1357 488
rect -933 -488 -899 488
rect -475 -488 -441 488
rect -17 -488 17 488
rect 441 -488 475 488
rect 899 -488 933 488
rect 1357 -488 1391 488
rect 1815 -488 1849 488
rect 2273 -488 2307 488
rect 2731 -488 2765 488
rect 3189 -488 3223 488
rect 3647 -488 3681 488
rect 4105 -488 4139 488
rect 4563 -488 4597 488
rect -4425 -581 -4277 -547
rect -3967 -581 -3819 -547
rect -3509 -581 -3361 -547
rect -3051 -581 -2903 -547
rect -2593 -581 -2445 -547
rect -2135 -581 -1987 -547
rect -1677 -581 -1529 -547
rect -1219 -581 -1071 -547
rect -761 -581 -613 -547
rect -303 -581 -155 -547
rect 155 -581 303 -547
rect 613 -581 761 -547
rect 1071 -581 1219 -547
rect 1529 -581 1677 -547
rect 1987 -581 2135 -547
rect 2445 -581 2593 -547
rect 2903 -581 3051 -547
rect 3361 -581 3509 -547
rect 3819 -581 3967 -547
rect 4277 -581 4425 -547
<< metal1 >>
rect -4437 581 -4265 587
rect -4437 547 -4425 581
rect -4277 547 -4265 581
rect -4437 541 -4265 547
rect -3979 581 -3807 587
rect -3979 547 -3967 581
rect -3819 547 -3807 581
rect -3979 541 -3807 547
rect -3521 581 -3349 587
rect -3521 547 -3509 581
rect -3361 547 -3349 581
rect -3521 541 -3349 547
rect -3063 581 -2891 587
rect -3063 547 -3051 581
rect -2903 547 -2891 581
rect -3063 541 -2891 547
rect -2605 581 -2433 587
rect -2605 547 -2593 581
rect -2445 547 -2433 581
rect -2605 541 -2433 547
rect -2147 581 -1975 587
rect -2147 547 -2135 581
rect -1987 547 -1975 581
rect -2147 541 -1975 547
rect -1689 581 -1517 587
rect -1689 547 -1677 581
rect -1529 547 -1517 581
rect -1689 541 -1517 547
rect -1231 581 -1059 587
rect -1231 547 -1219 581
rect -1071 547 -1059 581
rect -1231 541 -1059 547
rect -773 581 -601 587
rect -773 547 -761 581
rect -613 547 -601 581
rect -773 541 -601 547
rect -315 581 -143 587
rect -315 547 -303 581
rect -155 547 -143 581
rect -315 541 -143 547
rect 143 581 315 587
rect 143 547 155 581
rect 303 547 315 581
rect 143 541 315 547
rect 601 581 773 587
rect 601 547 613 581
rect 761 547 773 581
rect 601 541 773 547
rect 1059 581 1231 587
rect 1059 547 1071 581
rect 1219 547 1231 581
rect 1059 541 1231 547
rect 1517 581 1689 587
rect 1517 547 1529 581
rect 1677 547 1689 581
rect 1517 541 1689 547
rect 1975 581 2147 587
rect 1975 547 1987 581
rect 2135 547 2147 581
rect 1975 541 2147 547
rect 2433 581 2605 587
rect 2433 547 2445 581
rect 2593 547 2605 581
rect 2433 541 2605 547
rect 2891 581 3063 587
rect 2891 547 2903 581
rect 3051 547 3063 581
rect 2891 541 3063 547
rect 3349 581 3521 587
rect 3349 547 3361 581
rect 3509 547 3521 581
rect 3349 541 3521 547
rect 3807 581 3979 587
rect 3807 547 3819 581
rect 3967 547 3979 581
rect 3807 541 3979 547
rect 4265 581 4437 587
rect 4265 547 4277 581
rect 4425 547 4437 581
rect 4265 541 4437 547
rect -4603 488 -4557 500
rect -4603 -488 -4597 488
rect -4563 -488 -4557 488
rect -4603 -500 -4557 -488
rect -4145 488 -4099 500
rect -4145 -488 -4139 488
rect -4105 -488 -4099 488
rect -4145 -500 -4099 -488
rect -3687 488 -3641 500
rect -3687 -488 -3681 488
rect -3647 -488 -3641 488
rect -3687 -500 -3641 -488
rect -3229 488 -3183 500
rect -3229 -488 -3223 488
rect -3189 -488 -3183 488
rect -3229 -500 -3183 -488
rect -2771 488 -2725 500
rect -2771 -488 -2765 488
rect -2731 -488 -2725 488
rect -2771 -500 -2725 -488
rect -2313 488 -2267 500
rect -2313 -488 -2307 488
rect -2273 -488 -2267 488
rect -2313 -500 -2267 -488
rect -1855 488 -1809 500
rect -1855 -488 -1849 488
rect -1815 -488 -1809 488
rect -1855 -500 -1809 -488
rect -1397 488 -1351 500
rect -1397 -488 -1391 488
rect -1357 -488 -1351 488
rect -1397 -500 -1351 -488
rect -939 488 -893 500
rect -939 -488 -933 488
rect -899 -488 -893 488
rect -939 -500 -893 -488
rect -481 488 -435 500
rect -481 -488 -475 488
rect -441 -488 -435 488
rect -481 -500 -435 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 435 488 481 500
rect 435 -488 441 488
rect 475 -488 481 488
rect 435 -500 481 -488
rect 893 488 939 500
rect 893 -488 899 488
rect 933 -488 939 488
rect 893 -500 939 -488
rect 1351 488 1397 500
rect 1351 -488 1357 488
rect 1391 -488 1397 488
rect 1351 -500 1397 -488
rect 1809 488 1855 500
rect 1809 -488 1815 488
rect 1849 -488 1855 488
rect 1809 -500 1855 -488
rect 2267 488 2313 500
rect 2267 -488 2273 488
rect 2307 -488 2313 488
rect 2267 -500 2313 -488
rect 2725 488 2771 500
rect 2725 -488 2731 488
rect 2765 -488 2771 488
rect 2725 -500 2771 -488
rect 3183 488 3229 500
rect 3183 -488 3189 488
rect 3223 -488 3229 488
rect 3183 -500 3229 -488
rect 3641 488 3687 500
rect 3641 -488 3647 488
rect 3681 -488 3687 488
rect 3641 -500 3687 -488
rect 4099 488 4145 500
rect 4099 -488 4105 488
rect 4139 -488 4145 488
rect 4099 -500 4145 -488
rect 4557 488 4603 500
rect 4557 -488 4563 488
rect 4597 -488 4603 488
rect 4557 -500 4603 -488
rect -4437 -547 -4265 -541
rect -4437 -581 -4425 -547
rect -4277 -581 -4265 -547
rect -4437 -587 -4265 -581
rect -3979 -547 -3807 -541
rect -3979 -581 -3967 -547
rect -3819 -581 -3807 -547
rect -3979 -587 -3807 -581
rect -3521 -547 -3349 -541
rect -3521 -581 -3509 -547
rect -3361 -581 -3349 -547
rect -3521 -587 -3349 -581
rect -3063 -547 -2891 -541
rect -3063 -581 -3051 -547
rect -2903 -581 -2891 -547
rect -3063 -587 -2891 -581
rect -2605 -547 -2433 -541
rect -2605 -581 -2593 -547
rect -2445 -581 -2433 -547
rect -2605 -587 -2433 -581
rect -2147 -547 -1975 -541
rect -2147 -581 -2135 -547
rect -1987 -581 -1975 -547
rect -2147 -587 -1975 -581
rect -1689 -547 -1517 -541
rect -1689 -581 -1677 -547
rect -1529 -581 -1517 -547
rect -1689 -587 -1517 -581
rect -1231 -547 -1059 -541
rect -1231 -581 -1219 -547
rect -1071 -581 -1059 -547
rect -1231 -587 -1059 -581
rect -773 -547 -601 -541
rect -773 -581 -761 -547
rect -613 -581 -601 -547
rect -773 -587 -601 -581
rect -315 -547 -143 -541
rect -315 -581 -303 -547
rect -155 -581 -143 -547
rect -315 -587 -143 -581
rect 143 -547 315 -541
rect 143 -581 155 -547
rect 303 -581 315 -547
rect 143 -587 315 -581
rect 601 -547 773 -541
rect 601 -581 613 -547
rect 761 -581 773 -547
rect 601 -587 773 -581
rect 1059 -547 1231 -541
rect 1059 -581 1071 -547
rect 1219 -581 1231 -547
rect 1059 -587 1231 -581
rect 1517 -547 1689 -541
rect 1517 -581 1529 -547
rect 1677 -581 1689 -547
rect 1517 -587 1689 -581
rect 1975 -547 2147 -541
rect 1975 -581 1987 -547
rect 2135 -581 2147 -547
rect 1975 -587 2147 -581
rect 2433 -547 2605 -541
rect 2433 -581 2445 -547
rect 2593 -581 2605 -547
rect 2433 -587 2605 -581
rect 2891 -547 3063 -541
rect 2891 -581 2903 -547
rect 3051 -581 3063 -547
rect 2891 -587 3063 -581
rect 3349 -547 3521 -541
rect 3349 -581 3361 -547
rect 3509 -581 3521 -547
rect 3349 -587 3521 -581
rect 3807 -547 3979 -541
rect 3807 -581 3819 -547
rect 3967 -581 3979 -547
rect 3807 -587 3979 -581
rect 4265 -547 4437 -541
rect 4265 -581 4277 -547
rect 4425 -581 4437 -547
rect 4265 -587 4437 -581
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string parameters w 5 l 2 m 1 nf 20 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 40 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
