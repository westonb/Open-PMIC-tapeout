magic
tech sky130A
magscale 1 2
timestamp 1622500023
<< nwell >>
rect -2600 3700 8900 9000
<< pwell >>
rect -2600 0 8900 3600
rect 9100 0 11000 7200
<< mvpsubdiff >>
rect 9166 7122 10934 7134
rect 9166 6962 9400 7122
rect 10700 6962 10934 7122
rect 9166 6950 10934 6962
rect 9166 6900 9350 6950
rect -2534 3522 8834 3534
rect -2534 3362 -2300 3522
rect 8600 3362 8834 3522
rect -2534 3350 8834 3362
rect -2534 3300 -2350 3350
rect -2534 300 -2522 3300
rect -2362 300 -2350 3300
rect -2534 250 -2350 300
rect 8650 3300 8834 3350
rect 8650 300 8662 3300
rect 8822 300 8834 3300
rect 8650 250 8834 300
rect -2534 238 8834 250
rect -2534 78 -2300 238
rect 8600 78 8834 238
rect -2534 66 8834 78
rect 9166 300 9178 6900
rect 9338 300 9350 6900
rect 9166 250 9350 300
rect 10750 6900 10934 6950
rect 10750 300 10762 6900
rect 10922 300 10934 6900
rect 10750 250 10934 300
rect 9166 238 10934 250
rect 9166 78 9400 238
rect 10700 78 10934 238
rect 9166 66 10934 78
<< mvnsubdiff >>
rect -2534 8922 8834 8934
rect -2534 8762 -2300 8922
rect 8600 8762 8834 8922
rect -2534 8750 8834 8762
rect -2534 8700 -2350 8750
rect -2534 4000 -2522 8700
rect -2362 4000 -2350 8700
rect -2534 3950 -2350 4000
rect 8650 8700 8834 8750
rect 8650 4000 8662 8700
rect 8822 4000 8834 8700
rect 8650 3950 8834 4000
rect -2534 3938 8834 3950
rect -2534 3778 -2300 3938
rect 8600 3778 8834 3938
rect -2534 3766 8834 3778
<< mvpsubdiffcont >>
rect 9400 6962 10700 7122
rect -2300 3362 8600 3522
rect -2522 300 -2362 3300
rect 8662 300 8822 3300
rect -2300 78 8600 238
rect 9178 300 9338 6900
rect 10762 300 10922 6900
rect 9400 78 10700 238
<< mvnsubdiffcont >>
rect -2300 8762 8600 8922
rect -2522 4000 -2362 8700
rect 8662 4000 8822 8700
rect -2300 3778 8600 3938
<< locali >>
rect -2522 8700 -2362 8922
rect 8662 8700 8822 8922
rect -881 6853 -847 6896
rect 35 6853 69 6896
rect 951 6853 985 6896
rect 4615 6853 4649 6896
rect 5531 6853 5565 6896
rect 6447 6853 6481 6896
rect -1219 6785 1495 6853
rect 1815 6785 3785 6853
rect 4105 6785 6819 6853
rect -1219 6453 6819 6785
rect -1291 5747 5291 6247
rect 1983 5704 2017 5747
rect 6983 4653 7017 4696
rect 6289 4453 7745 4653
rect -2522 3778 -2362 4000
rect 8662 3778 8822 4000
rect 9178 6900 9338 7122
rect -2522 3300 -2362 3522
rect 8662 3300 8822 3522
rect 2331 2638 2979 2713
rect 1815 2613 3237 2638
rect 1815 2538 2463 2613
rect 2847 2538 3237 2613
rect 3363 2538 4785 2638
rect 6455 2538 6513 2572
rect 1993 2504 2027 2538
rect 3025 2504 3059 2538
rect 3541 2504 3575 2538
rect 4573 2504 4607 2538
rect 5615 2466 5677 2538
rect 5773 2466 5835 2538
rect 5869 2466 5931 2538
rect 6027 2466 6089 2538
rect 6247 2466 6309 2538
rect 6405 2504 6563 2538
rect 6405 2466 6467 2504
rect 6501 2466 6563 2504
rect 6659 2466 6721 2538
rect 6879 2466 6941 2538
rect 7037 2466 7099 2538
rect 7133 2466 7195 2538
rect 7291 2466 7353 2538
rect 7511 2466 7573 2538
rect 7669 2466 7731 2538
rect 7765 2466 7827 2538
rect 7923 2466 7985 2538
rect 5361 1462 5395 1496
rect 8205 1462 8239 1496
rect 5361 1428 5507 1462
rect 8093 1428 8239 1462
rect -2522 78 -2362 300
rect 8662 78 8822 300
rect 9178 78 9338 300
rect 10762 6900 10922 7122
rect 10762 78 10922 300
<< viali >>
rect -2362 8762 -2300 8922
rect -2300 8762 8600 8922
rect 8600 8762 8662 8922
rect -2522 4179 -2362 8521
rect 8662 4179 8822 8521
rect -2362 3778 -2300 3938
rect -2300 3778 8600 3938
rect 8600 3778 8662 3938
rect 9338 6962 9400 7122
rect 9400 6962 10700 7122
rect 10700 6962 10762 7122
rect -2362 3362 -2300 3522
rect -2300 3362 8600 3522
rect 8600 3362 8662 3522
rect -2522 394 -2362 3206
rect 8662 394 8822 3206
rect -2362 78 -2300 238
rect -2300 78 8600 238
rect 8600 78 8662 238
rect 9178 574 9338 6626
rect 10762 574 10922 6626
rect 9338 78 9400 238
rect 9400 78 10700 238
rect 10700 78 10762 238
<< metal1 >>
rect -2528 8922 8828 8928
rect -2528 8762 -2362 8922
rect 8662 8762 8828 8922
rect -2528 8756 8828 8762
rect -2528 8521 -2356 8756
rect -2528 4179 -2522 8521
rect -2362 8456 -2356 8521
rect -1756 8456 8056 8756
rect 8656 8521 8828 8756
rect 8656 8456 8662 8521
rect -2362 8380 8662 8456
rect -2362 6340 -1937 8380
rect -1803 8140 7403 8380
rect -1803 7987 -1757 8140
rect -1803 7941 -1465 7987
rect -1803 7900 -1757 7941
rect -1345 7900 -1299 8140
rect -429 7900 -383 8140
rect 487 7900 533 8140
rect 1403 7987 1449 8140
rect 3693 7987 3739 8140
rect 4151 7987 4197 8140
rect 1403 7941 1741 7987
rect 3693 7941 4197 7987
rect 1403 7900 1449 7941
rect 3693 7900 3739 7941
rect 4151 7900 4197 7941
rect 5067 7900 5113 8140
rect 5983 7900 6029 8140
rect 6899 7900 6945 8140
rect 7357 7987 7403 8140
rect 7065 7941 7403 7987
rect 7357 7900 7403 7941
rect -887 6660 -841 6900
rect 29 6660 75 6900
rect 945 6660 991 6900
rect 1861 6806 1907 6900
rect 1848 6754 1858 6806
rect 1910 6754 1920 6806
rect 4609 6660 4655 6900
rect 5525 6660 5571 6900
rect 6441 6660 6487 6900
rect -887 6638 6487 6660
rect -887 6586 2767 6638
rect 2819 6586 6487 6638
rect -887 6560 6487 6586
rect 7804 6340 8662 8380
rect -2362 5940 8662 6340
rect -2362 4179 -2356 5940
rect -1635 5787 -1589 5940
rect -1377 5787 -1331 5940
rect -1635 5741 -1331 5787
rect -1635 5700 -1589 5741
rect -1377 5700 -1331 5741
rect -861 5700 -815 5940
rect -345 5700 -299 5940
rect 171 5700 217 5940
rect 687 5700 733 5940
rect 1203 5700 1249 5940
rect 1719 5700 1765 5940
rect 1964 5794 1974 5846
rect 2026 5794 2036 5846
rect 1964 5787 2036 5794
rect 1825 5741 2175 5787
rect 1977 5700 2023 5741
rect 2235 5700 2281 5940
rect 2751 5700 2797 5940
rect 3267 5700 3313 5940
rect 3783 5700 3829 5940
rect 4299 5700 4345 5940
rect 4815 5700 4861 5940
rect 5331 5787 5377 5940
rect 5589 5787 5635 5940
rect 5331 5741 5635 5787
rect 5331 5700 5377 5741
rect 5589 5700 5635 5741
rect 5945 5787 5991 5940
rect 6203 5787 6249 5940
rect 5945 5741 6249 5787
rect 5945 5700 5991 5741
rect 6203 5700 6249 5741
rect 6719 5700 6765 5940
rect 7235 5700 7281 5940
rect 7751 5787 7797 5940
rect 8009 5787 8055 5940
rect 7751 5741 8055 5787
rect 7751 5700 7797 5741
rect 8009 5700 8055 5741
rect -1119 4460 -1073 4700
rect -603 4460 -557 4700
rect -87 4606 -41 4700
rect -100 4554 -90 4606
rect -38 4554 -28 4606
rect 429 4460 475 4700
rect 945 4606 991 4700
rect 932 4554 942 4606
rect 994 4554 1004 4606
rect 1461 4460 1507 4700
rect 2493 4460 2539 4700
rect 3009 4606 3055 4700
rect 2996 4554 3006 4606
rect 3058 4554 3068 4606
rect 3525 4460 3571 4700
rect 4041 4606 4087 4700
rect 4028 4554 4038 4606
rect 4090 4554 4100 4606
rect 4557 4460 4603 4700
rect 5073 4460 5119 4700
rect -1119 4415 5119 4460
rect -1119 4220 1907 4415
rect 1897 4215 1907 4220
rect 2107 4220 5119 4415
rect 5501 4459 5601 4465
rect 6461 4460 6507 4700
rect 6977 4659 7023 4700
rect 6825 4613 7175 4659
rect 6964 4606 7036 4613
rect 6964 4554 6974 4606
rect 7026 4554 7036 4606
rect 7493 4460 7539 4700
rect 6461 4459 7539 4460
rect 5601 4432 7539 4459
rect 5601 4380 7116 4432
rect 7168 4380 7539 4432
rect 5601 4359 7539 4380
rect 5501 4353 5601 4359
rect 2107 4215 2117 4220
rect -2528 3944 -2356 4179
rect 8656 4179 8662 5940
rect 8822 4179 8828 8521
rect 8656 3944 8828 4179
rect -2528 3938 8828 3944
rect -2528 3778 -2362 3938
rect 8662 3778 8828 3938
rect -2528 3772 8828 3778
rect 9172 7122 10928 7128
rect 9172 6962 9338 7122
rect 10762 6962 10928 7122
rect 9172 6956 10928 6962
rect 9172 6626 9344 6956
rect -2528 3522 8828 3528
rect -2528 3362 -2362 3522
rect 8662 3362 8828 3522
rect -2528 3356 8828 3362
rect -2528 3206 -2356 3356
rect -2737 1772 -2731 1852
rect -2651 1772 -2645 1852
rect -2731 678 -2651 1772
rect -2731 592 -2651 598
rect -2528 394 -2522 3206
rect -2362 610 -2356 3206
rect 8656 3206 8828 3356
rect 109 2940 115 2948
rect -2051 2919 115 2940
rect -2051 2827 -643 2919
rect -551 2827 115 2919
rect -2051 2748 115 2827
rect 315 2940 321 2948
rect 315 2748 397 2940
rect -2051 2740 397 2748
rect -2051 1560 -1851 2740
rect -1197 2500 -1151 2740
rect -681 2500 -635 2740
rect -436 2594 -426 2646
rect -374 2594 -364 2646
rect -423 2500 -377 2594
rect -165 2500 -119 2740
rect 351 2500 397 2740
rect 1081 2882 3915 2962
rect -2051 1354 -1851 1360
rect -1713 1468 -1667 1500
rect -1455 1468 -1409 1500
rect -1713 1422 -1409 1468
rect -1713 1260 -1667 1422
rect -1455 1260 -1409 1422
rect -1349 1428 -999 1468
rect -1349 1376 -1200 1428
rect -1148 1376 -999 1428
rect -1349 1368 -999 1376
rect -939 1260 -893 1500
rect -833 1428 33 1468
rect -833 1376 -427 1428
rect -375 1376 33 1428
rect -833 1368 33 1376
rect 93 1260 139 1500
rect 609 1468 655 1500
rect 867 1468 913 1500
rect 199 1428 549 1468
rect 199 1376 348 1428
rect 400 1376 549 1428
rect 199 1368 549 1376
rect 609 1422 913 1468
rect 609 1260 655 1422
rect 867 1260 913 1422
rect -1713 610 913 1260
rect 1081 955 1161 2882
rect 3835 2820 3915 2882
rect 1081 869 1161 875
rect 1243 2740 3065 2820
rect 1243 768 1323 2740
rect 1987 2500 2033 2740
rect 2490 2594 2500 2646
rect 2552 2594 2562 2646
rect 2503 2500 2549 2594
rect 3019 2500 3065 2740
rect 3535 2740 4613 2820
rect 3535 2500 3581 2740
rect 4038 2594 4048 2646
rect 4100 2594 4110 2646
rect 4051 2500 4097 2594
rect 4567 2500 4613 2740
rect 5671 2740 7929 2820
rect 5671 2500 5717 2740
rect 5816 2594 5826 2646
rect 5878 2594 5888 2646
rect 5829 2500 5875 2594
rect 5987 2500 6033 2740
rect 6303 2500 6349 2740
rect 6448 2594 6458 2646
rect 6510 2594 6520 2646
rect 6461 2500 6507 2594
rect 6619 2500 6665 2740
rect 6935 2500 6981 2740
rect 7080 2594 7090 2646
rect 7142 2594 7152 2646
rect 7093 2500 7139 2594
rect 7251 2500 7297 2740
rect 7567 2500 7613 2740
rect 7712 2594 7722 2646
rect 7774 2594 7784 2646
rect 7725 2500 7771 2594
rect 7883 2500 7929 2740
rect 1471 1468 1517 1500
rect 1729 1468 1775 1500
rect 1471 1422 1775 1468
rect 1471 1260 1517 1422
rect 1729 1260 1775 1422
rect 2245 1260 2291 1500
rect 2761 1468 2807 1500
rect 2609 1422 2807 1468
rect 2761 1260 2807 1422
rect 3277 1260 3323 1500
rect 3793 1260 3839 1500
rect 4309 1260 4355 1500
rect 4825 1468 4871 1500
rect 5083 1468 5129 1500
rect 4825 1422 5129 1468
rect 4825 1260 4871 1422
rect 5083 1260 5129 1422
rect 1096 767 1323 768
rect 1038 687 1044 767
rect 1124 688 1323 767
rect 1124 687 1207 688
rect 1472 610 5129 1260
rect 5355 1260 5401 1500
rect 5513 1260 5559 1500
rect 6145 1260 6191 1500
rect 6777 1260 6823 1500
rect 7409 1260 7455 1500
rect 8041 1260 8087 1500
rect 8199 1260 8245 1500
rect 5355 610 8245 1260
rect 8656 610 8662 3206
rect -2362 544 8662 610
rect -2362 394 -2356 544
rect -2528 244 -2356 394
rect -1756 244 8056 544
rect 8656 394 8662 544
rect 8822 394 8828 3206
rect 8656 244 8828 394
rect -2528 238 8828 244
rect -2528 78 -2362 238
rect 8662 78 8828 238
rect -2528 72 8828 78
rect 9172 574 9178 6626
rect 9338 574 9344 6626
rect 10756 6626 10928 6956
rect 9921 5819 10021 5825
rect 9921 5713 10021 5719
rect 9172 244 9344 574
rect 9839 544 10188 1489
rect 10756 574 10762 6626
rect 10922 574 10928 6626
rect 9944 244 10156 544
rect 10756 244 10928 574
rect 9172 238 10928 244
rect 9172 78 9338 238
rect 10762 78 10928 238
rect 9172 72 10928 78
<< via1 >>
rect -2356 8456 -1756 8756
rect 8056 8456 8656 8756
rect 1858 6754 1910 6806
rect 2767 6586 2819 6638
rect 1974 5794 2026 5846
rect -90 4554 -38 4606
rect 942 4554 994 4606
rect 3006 4554 3058 4606
rect 4038 4554 4090 4606
rect 1907 4215 2107 4415
rect 6974 4554 7026 4606
rect 5501 4359 5601 4459
rect 7116 4380 7168 4432
rect -2731 1772 -2651 1852
rect -2731 598 -2651 678
rect -643 2827 -551 2919
rect 115 2748 315 2948
rect -426 2594 -374 2646
rect -2051 1360 -1851 1560
rect -1200 1376 -1148 1428
rect -427 1376 -375 1428
rect 348 1376 400 1428
rect 1081 875 1161 955
rect 2500 2594 2552 2646
rect 4048 2594 4100 2646
rect 5826 2594 5878 2646
rect 6458 2594 6510 2646
rect 7090 2594 7142 2646
rect 7722 2594 7774 2646
rect 1044 687 1124 767
rect -2356 244 -1756 544
rect 8056 244 8656 544
rect 9921 5719 10021 5819
rect 9344 244 9944 544
rect 10156 244 10756 544
<< metal2 >>
rect -2356 8756 -1756 8766
rect -2356 8446 -1756 8456
rect 8056 8756 8656 8766
rect 8056 8446 8656 8456
rect 1844 6806 1924 6816
rect 1844 6754 1858 6806
rect 1910 6754 1924 6806
rect 1844 6596 1924 6754
rect -2250 6516 1924 6596
rect 2753 6638 2833 6648
rect 2753 6586 2767 6638
rect 2819 6586 2833 6638
rect -2250 4104 -2170 6516
rect 2753 6514 2833 6586
rect 2753 6434 5791 6514
rect -2021 5905 1835 5977
rect -2021 4116 -1949 5905
rect 1763 5856 1835 5905
rect 1763 5846 2026 5856
rect 1763 5794 1974 5846
rect 1763 5784 2026 5794
rect -90 4606 -38 4616
rect 942 4606 994 4616
rect 3006 4606 3058 4616
rect 4038 4606 4090 4616
rect -38 4554 942 4606
rect 994 4554 3006 4606
rect 3058 4554 4038 4606
rect 4090 4554 4261 4606
rect -90 4506 4261 4554
rect 4161 4459 4261 4506
rect 1907 4415 2107 4425
rect 4161 4359 5501 4459
rect 5601 4359 5607 4459
rect -2731 4024 -2170 4104
rect -2030 4044 -2021 4116
rect -1949 4044 -1940 4116
rect -2731 3040 -2651 4024
rect 1907 3200 2107 4215
rect 5711 3331 5791 6434
rect 8442 5719 9921 5819
rect 10021 5719 10027 5819
rect -2731 2960 -360 3040
rect -2731 2005 -2651 2960
rect -643 2919 -551 2925
rect -2839 1995 -2651 2005
rect -2750 1923 -2651 1995
rect -2839 1913 -2651 1923
rect -2731 1852 -2651 1913
rect -2731 1766 -2651 1772
rect -2510 2827 -643 2919
rect -2510 1694 -2418 2827
rect -643 2821 -551 2827
rect -440 2646 -360 2960
rect 115 3000 2107 3200
rect 3799 3251 5791 3331
rect 6955 4606 7055 4635
rect 6955 4554 6974 4606
rect 7026 4554 7055 4606
rect 3799 3090 3879 3251
rect 6955 3121 7055 4554
rect 8442 4460 8542 5719
rect 7116 4432 8542 4460
rect 7168 4380 8542 4432
rect 7116 4360 8542 4380
rect 2489 3010 3879 3090
rect 4024 3021 7055 3121
rect 115 2948 315 3000
rect 115 2742 315 2748
rect -440 2594 -426 2646
rect -374 2594 -360 2646
rect -440 2584 -360 2594
rect -3100 1689 -2418 1694
rect -3104 1619 -3095 1689
rect -3025 1619 -2418 1689
rect -3100 1614 -2418 1619
rect -2510 1370 -2418 1614
rect -2597 1360 -2357 1370
rect -2057 1360 -2051 1560
rect -1851 1360 -1845 1560
rect -1200 1428 400 1438
rect -1148 1376 -427 1428
rect -375 1376 348 1428
rect -1200 1366 400 1376
rect -4584 1023 -4575 1223
rect -4375 1038 -4003 1223
rect -2597 1110 -2357 1120
rect -2051 1038 -1851 1360
rect -711 1166 -639 1366
rect -711 1085 -639 1094
rect -4375 1023 -1851 1038
rect -4583 838 -1851 1023
rect -1620 875 -1611 955
rect -1531 875 1081 955
rect 1161 875 1167 955
rect 1044 767 1124 773
rect -6808 652 -6736 657
rect -6812 590 -6803 652
rect -6741 590 -6732 652
rect -2737 598 -2731 678
rect -2651 598 -2645 678
rect -7014 434 -6944 438
rect -7019 429 -6939 434
rect -7019 359 -7014 429
rect -6944 359 -6939 429
rect -7019 -5799 -6939 359
rect -10321 -5879 -10312 -5799
rect -10232 -5879 -6939 -5799
rect -6808 -6045 -6736 590
rect -2731 556 -2651 598
rect -2740 476 -2731 556
rect -2651 476 -2642 556
rect -2374 544 -1734 568
rect -6315 376 -6235 381
rect -6319 306 -6310 376
rect -6240 306 -6231 376
rect -10400 -6117 -10391 -6045
rect -10319 -6117 -6736 -6045
rect -6551 89 -6471 99
rect -6551 -6359 -6471 9
rect -10464 -6439 -10455 -6359
rect -10375 -6439 -6471 -6359
rect -6315 -6532 -6235 306
rect -2374 244 -2356 544
rect -1756 244 -1734 544
rect -2374 230 -1734 244
rect 1044 84 1124 687
rect 1044 14 1049 84
rect 1119 14 1124 84
rect 1044 9 1124 14
rect 1049 5 1119 9
rect -6139 -563 -6049 -559
rect -6144 -568 -6044 -563
rect -6144 -658 -6139 -568
rect -6049 -658 -6044 -568
rect -6144 -3727 -6044 -658
rect -6144 -3797 -6128 -3727
rect -6058 -3797 -6044 -3727
rect -6144 -4772 -6044 -3797
rect -6144 -4881 -6044 -4872
rect -6324 -6612 -6315 -6532
rect -6235 -6612 -6226 -6532
rect 1288 -6553 1348 3000
rect 2489 2646 2569 3010
rect 2489 2594 2500 2646
rect 2552 2594 2569 2646
rect 2489 2581 2569 2594
rect 4024 2646 4124 3021
rect 4024 2594 4048 2646
rect 4100 2594 4124 2646
rect 4024 2584 4124 2594
rect 5211 2646 7774 2684
rect 5211 2594 5826 2646
rect 5878 2594 6458 2646
rect 6510 2594 7090 2646
rect 7142 2594 7722 2646
rect 5211 2584 7774 2594
rect 5211 1068 5311 2584
rect 2500 968 5311 1068
rect 2507 -563 2607 968
rect 8948 805 9048 5719
rect 2755 800 2855 805
rect 2751 710 2760 800
rect 2850 710 2859 800
rect 2507 -672 2607 -663
rect 2755 -4814 2855 710
rect 8414 705 8423 805
rect 8523 705 9048 805
rect 8056 544 8656 554
rect 8056 234 8656 244
rect 9344 544 9944 554
rect 9344 234 9944 244
rect 10156 544 10756 554
rect 10156 234 10756 244
rect 2755 -4870 2783 -4814
rect 2839 -4870 2855 -4814
rect 2755 -4889 2855 -4870
rect 1281 -6609 1290 -6553
rect 1346 -6609 1355 -6553
rect 1288 -6611 1348 -6609
<< via2 >>
rect -2356 8456 -1756 8756
rect 8056 8456 8656 8756
rect -2021 4044 -1949 4116
rect -2839 1923 -2750 1995
rect -3095 1619 -3025 1689
rect -4575 1023 -4375 1223
rect -2597 1120 -2357 1360
rect -711 1094 -639 1166
rect -1611 875 -1531 955
rect -6803 590 -6741 652
rect -7014 359 -6944 429
rect -10312 -5879 -10232 -5799
rect -2731 476 -2651 556
rect -6310 306 -6240 376
rect -10391 -6117 -10319 -6045
rect -6551 9 -6471 89
rect -10455 -6439 -10375 -6359
rect -2356 244 -1756 544
rect 1049 14 1119 84
rect -6139 -658 -6049 -568
rect -6128 -3797 -6058 -3727
rect -6144 -4872 -6044 -4772
rect -6315 -6612 -6235 -6532
rect 2760 710 2850 800
rect 2507 -663 2607 -563
rect 8423 705 8523 805
rect 8056 244 8656 544
rect 9344 244 9944 544
rect 10156 244 10756 544
rect 2783 -4870 2839 -4814
rect 1290 -6609 1346 -6553
<< metal3 >>
rect -2366 8756 -1746 8761
rect -2366 8456 -2356 8756
rect -1756 8456 -1746 8756
rect -2366 8451 -1746 8456
rect 8046 8756 8666 8761
rect 8046 8456 8056 8756
rect 8656 8456 8666 8756
rect 8046 8451 8666 8456
rect -9700 2097 -3100 8000
rect -2026 4116 -1944 4121
rect -2026 4044 -2021 4116
rect -1949 4044 -1944 4116
rect -2026 4039 -1944 4044
rect -2021 3705 -1949 4039
rect -2265 3633 -1949 3705
rect -9700 1800 -3020 2097
rect -2915 1840 -2905 2055
rect -2668 1840 -2658 2055
rect -3100 1689 -3020 1800
rect -3100 1619 -3095 1689
rect -3025 1619 -3020 1689
rect -3100 1614 -3020 1619
rect -2607 1360 -2347 1365
rect -10318 1223 -4370 1228
rect -10318 1023 -4575 1223
rect -4375 1023 -4370 1223
rect -2607 1120 -2597 1360
rect -2357 1120 -2347 1360
rect -2607 1115 -2347 1120
rect -10318 828 -4370 1023
rect -2265 1003 -2193 3633
rect -716 1166 -634 1171
rect -716 1094 -711 1166
rect -639 1094 -634 1166
rect -716 1089 -634 1094
rect -4262 931 -2193 1003
rect -1616 955 -1526 960
rect -4262 748 -4190 931
rect -2032 875 -1611 955
rect -1531 875 -1526 955
rect -2032 869 -1952 875
rect -1616 870 -1526 875
rect -6808 676 -4190 748
rect -4067 789 -1952 869
rect -6808 652 -6736 676
rect -6808 590 -6803 652
rect -6741 590 -6736 652
rect -6808 585 -6736 590
rect -4067 579 -3982 789
rect -6510 499 -3982 579
rect -2736 556 -2646 561
rect -6510 434 -6430 499
rect -7019 429 -6430 434
rect -7019 359 -7014 429
rect -6944 359 -6430 429
rect -3756 476 -2731 556
rect -2651 476 -2646 556
rect -3756 381 -3676 476
rect -2736 471 -2646 476
rect -2366 544 -1746 549
rect -7019 354 -6430 359
rect -6315 376 -3676 381
rect -6315 306 -6310 376
rect -6240 306 -3676 376
rect -6315 301 -3676 306
rect -2366 244 -2356 544
rect -1756 244 -1746 544
rect -711 356 -639 1089
rect 8418 805 8528 810
rect 2755 800 8423 805
rect 2755 710 2760 800
rect 2850 710 8423 800
rect 2755 705 8423 710
rect 8523 705 8528 805
rect 8418 700 8528 705
rect 8046 544 8666 549
rect -711 284 3542 356
rect -2366 239 -1746 244
rect -6556 89 -6466 94
rect -6556 9 -6551 89
rect -6471 84 1124 89
rect -6471 14 1049 84
rect 1119 14 1124 84
rect -6471 9 1124 14
rect 3470 40 3542 284
rect 8046 244 8056 544
rect 8656 244 8666 544
rect 8046 239 8666 244
rect 9334 544 9954 549
rect 9334 244 9344 544
rect 9944 244 9954 544
rect 9334 239 9954 244
rect 10146 544 10766 549
rect 10146 244 10156 544
rect 10756 244 10766 544
rect 10146 239 10766 244
rect -6556 4 -6466 9
rect 3470 -32 9110 40
rect 2502 -563 2612 -558
rect -6144 -568 2507 -563
rect -6144 -658 -6139 -568
rect -6049 -658 2507 -568
rect -6144 -663 2507 -658
rect 2607 -663 2612 -563
rect 2502 -668 2612 -663
rect 9038 -916 9110 -32
rect 9038 -988 11740 -916
rect -10496 -3727 -6053 -3722
rect -10496 -3797 -6128 -3727
rect -6058 -3797 -6053 -3727
rect -10496 -3802 -6053 -3797
rect 227 -4534 11792 -4474
rect -6149 -4772 -6039 -4767
rect -6149 -4872 -6144 -4772
rect -6044 -4872 -5561 -4772
rect -6149 -4877 -6039 -4872
rect 227 -5252 287 -4534
rect 2778 -4812 2844 -4809
rect 2778 -4814 3439 -4812
rect 2778 -4870 2783 -4814
rect 2839 -4870 3439 -4814
rect 2778 -4872 3439 -4870
rect 2778 -4875 2844 -4872
rect -326 -5312 287 -5252
rect 8663 -5326 11825 -5238
rect -10317 -5799 -10227 -5794
rect -10509 -5879 -10312 -5799
rect -10232 -5879 -10227 -5799
rect -10317 -5884 -10227 -5879
rect -10396 -6045 -10314 -6040
rect -10512 -6117 -10391 -6045
rect -10319 -6117 -10314 -6045
rect -10396 -6122 -10314 -6117
rect -10460 -6359 -10370 -6354
rect -10531 -6439 -10455 -6359
rect -10375 -6439 -10370 -6359
rect -10460 -6444 -10370 -6439
rect -6320 -6532 -6230 -6527
rect -6320 -6612 -6315 -6532
rect -6235 -6612 -5672 -6532
rect -6320 -6617 -6230 -6612
rect -5752 -6636 -5672 -6612
rect 1285 -6551 1351 -6548
rect 1285 -6553 3313 -6551
rect 1285 -6609 1290 -6553
rect 1346 -6609 3313 -6553
rect 1285 -6611 3313 -6609
rect 1285 -6614 1351 -6611
rect -5752 -6716 -5522 -6636
rect 3253 -6653 3313 -6611
rect 3253 -6713 3465 -6653
rect -10570 -6819 -6023 -6775
rect -10570 -6820 -5669 -6819
rect 2345 -6820 2904 -6780
rect -10570 -6880 -5573 -6820
rect 2345 -6880 3459 -6820
rect -10570 -6922 -6023 -6880
rect 2345 -6919 2904 -6880
rect -10586 -7410 -6250 -7271
rect -6389 -8235 -6250 -7410
rect 2345 -8192 2484 -6919
rect -6389 -8374 -4872 -8235
rect -5011 -8515 -4872 -8374
rect -1042 -8331 2484 -8192
rect -1042 -8515 -903 -8331
rect -5011 -8654 -903 -8515
<< via3 >>
rect -2356 8456 -1756 8756
rect 8056 8456 8656 8756
rect -2905 1995 -2668 2055
rect -2905 1923 -2839 1995
rect -2839 1923 -2750 1995
rect -2750 1923 -2668 1995
rect -2905 1840 -2668 1923
rect -2597 1120 -2357 1360
rect -2356 244 -1756 544
rect 8056 244 8656 544
rect 9344 244 9944 544
rect 10156 244 10756 544
<< mimcap >>
rect -9600 7850 -3200 7900
rect -9600 1950 -3550 7850
rect -3250 1950 -3200 7850
rect -9600 1900 -3200 1950
<< mimcapcontact >>
rect -3550 1950 -3250 7850
<< metal4 >>
rect -12000 8899 12000 9000
rect -12000 8299 -11817 8899
rect -10931 8756 12000 8899
rect -10931 8456 -2356 8756
rect -1756 8456 8056 8756
rect 8656 8456 12000 8756
rect -10931 8299 12000 8456
rect -12000 8200 12000 8299
rect -9700 7850 -3100 8000
rect -9700 1950 -3550 7850
rect -3250 2097 -3100 7850
rect -3250 2055 -2609 2097
rect -3250 1950 -2905 2055
rect -9700 1840 -2905 1950
rect -2668 1840 -2609 2055
rect -9700 1800 -2609 1840
rect -9700 1400 -3500 1800
rect -2598 1360 -2356 1361
rect -2598 1120 -2597 1360
rect -2357 1120 -2356 1360
rect -2598 1119 -2356 1120
rect -12000 544 12000 800
rect -12000 244 -2356 544
rect -1756 244 8056 544
rect 8656 244 9344 544
rect 9944 244 10156 544
rect 10756 244 12000 544
rect -12000 -800 12000 244
rect -12000 -8324 12000 -8200
rect -12000 -8924 -11844 -8324
rect -10958 -8924 12000 -8324
rect -12000 -9000 12000 -8924
<< via4 >>
rect -11817 8299 -10931 8899
rect -2597 1120 -2357 1360
rect -11844 -8924 -10958 -8324
<< mimcap2 >>
rect -9600 1850 -3600 7900
rect -9600 1550 -9550 1850
rect -3650 1550 -3600 1850
rect -9600 1500 -3600 1550
<< mimcap2contact >>
rect -9550 1550 -3650 1850
<< metal5 >>
rect -12000 8899 -10800 9000
rect -12000 8299 -11817 8899
rect -10931 8299 -10800 8899
rect -12000 -8324 -10800 8299
rect -9700 1850 -3500 8000
rect -9700 1550 -9550 1850
rect -3650 1550 -3500 1850
rect -9700 1400 -3500 1550
rect -3820 1360 -2317 1400
rect -3820 1120 -2597 1360
rect -2357 1120 -2317 1360
rect -3820 1080 -2317 1120
rect -12000 -8924 -11844 -8324
rect -10958 -8924 -10800 -8324
rect -12000 -9000 -10800 -8924
<< comment >>
rect 2772 6503 2818 6743
rect 1983 4407 2029 4647
rect -402 1118 -356 1358
rect 3283 1212 3329 1452
rect 6786 1093 6832 1333
use sky130_fd_pr__nfet_g5v0d10v5_V2YKKA  xm4
timestamp 1621758535
transform 1 0 -400 0 1 2000
box -1319 -588 1319 588
use comparator  comparator_1
timestamp 1621890638
transform 1 0 -3000 0 -1 -4500
box -3000 -4500 3000 4500
use comparator  comparator_0
timestamp 1621890638
transform 1 0 6000 0 -1 -4500
box -3000 -4500 3000 4500
use sky130_fd_pr__res_high_po_1p41_20um  sky130_fd_pr__res_high_po_1p41_20um_0
timestamp 1621741225
transform 1 0 10000 0 -1 3500
box -143 -2432 143 2432
use sky130_fd_pr__pfet_g5v0d10v5_QZEXLW  xm1
timestamp 1621838304
transform 1 0 2800 0 1 7400
box -4675 -600 4675 600
use sky130_fd_pr__pfet_g5v0d10v5_QVWX2D  xm2
timestamp 1621838304
transform 1 0 2000 0 1 5200
box -3707 -600 3707 600
use sky130_fd_pr__pfet_g5v0d10v5_ZBHAPX  xm3
timestamp 1621838304
transform 1 0 7000 0 1 5200
box -1127 -600 1127 600
use sky130_fd_pr__nfet_g5v0d10v5_DQEKNK  xm5
timestamp 1621838304
transform 1 0 3300 0 1 2000
box -1835 -588 1835 588
use sky130_fd_pr__nfet_g5v0d10v5_E8UHFU  xm6
timestamp 1621838304
transform 1 0 6800 0 1 2000
box -1451 -588 1451 588
<< labels >>
flabel metal4 -12000 8200 -12000 9000 3 FreeSans 480 0 0 0 vdd
port 11 e
flabel metal4 -12000 0 -12000 800 3 FreeSans 480 0 0 0 vss
port 12 e
flabel metal3 -10531 -6439 -10530 -6359 1 FreeSans 240 0 0 0 islope
port 7 n
flabel metal3 -10512 -6117 -10510 -6045 1 FreeSans 240 0 0 0 current_offset
port 3 n
flabel metal3 11823 -5326 11825 -5238 1 FreeSans 240 0 0 0 overcurrent
port 8 n
flabel metal3 11791 -4534 11792 -4474 1 FreeSans 240 0 0 0 cycle_end
port 4 n
flabel metal3 -10586 -7410 -10584 -7271 1 FreeSans 240 0 0 0 cmp_bias_2
port 2 n
flabel metal3 -10570 -6922 -10568 -6775 1 FreeSans 240 0 0 0 cmp_bias
port 1 n
flabel metal3 -10509 -5879 -10507 -5799 1 FreeSans 240 0 0 0 ioc
port 5 n
flabel metal3 -10496 -3802 -10494 -3722 1 FreeSans 240 0 0 0 vcomp
port 10 n
flabel metal3 -10318 828 -10314 1228 1 FreeSans 240 0 0 0 isense
port 6 n
flabel metal2 9786 5719 9788 5819 1 FreeSans 400 0 0 0 ioc_res
flabel metal2 -506 2960 -503 3040 1 FreeSans 400 0 0 0 imod
flabel metal2 2724 3010 2726 3090 1 FreeSans 400 0 0 0 islope_mirror
flabel metal3 11737 -988 11740 -916 1 FreeSans 400 0 0 0 timeout
port 9 n
<< properties >>
string FIXED_BBOX 9258 158 10842 7042
<< end >>
